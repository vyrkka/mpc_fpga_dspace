module motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config2_s (
        ap_clk,
        ap_rst,
        p_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [95:0] p_read;
output  [31:0] ap_return_0;
output  [31:0] ap_return_1;
output  [31:0] ap_return_2;
output  [31:0] ap_return_3;
output  [31:0] ap_return_4;
output  [31:0] ap_return_5;
output  [31:0] ap_return_6;
output  [31:0] ap_return_7;
output  [31:0] ap_return_8;
input   ap_ce;

reg[31:0] ap_return_0;
reg[31:0] ap_return_1;
reg[31:0] ap_return_2;
reg[31:0] ap_return_3;
reg[31:0] ap_return_4;
reg[31:0] ap_return_5;
reg[31:0] ap_return_6;
reg[31:0] ap_return_7;
reg[31:0] ap_return_8;

wire   [42:0] r_V_178_fu_254_p2;
reg   [42:0] r_V_178_reg_2283;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [43:0] r_V_179_fu_262_p2;
reg   [43:0] r_V_179_reg_2287;
wire   [56:0] r_V_180_fu_251_p2;
reg   [56:0] r_V_180_reg_2291;
wire   [43:0] r_V_181_fu_256_p2;
reg   [43:0] r_V_181_reg_2295;
wire   [46:0] r_V_182_fu_264_p2;
reg   [46:0] r_V_182_reg_2299;
wire   [42:0] r_V_183_fu_240_p2;
reg   [42:0] r_V_183_reg_2303;
wire   [42:0] r_V_184_fu_249_p2;
reg   [42:0] r_V_184_reg_2307;
wire   [53:0] r_V_185_fu_259_p2;
reg   [53:0] r_V_185_reg_2311;
wire   [53:0] r_V_186_fu_246_p2;
reg   [53:0] r_V_186_reg_2315;
wire   [40:0] r_V_187_fu_266_p2;
reg   [40:0] r_V_187_reg_2319;
wire   [42:0] r_V_188_fu_261_p2;
reg   [42:0] r_V_188_reg_2323;
wire   [44:0] r_V_189_fu_242_p2;
reg   [44:0] r_V_189_reg_2327;
wire   [42:0] r_V_190_fu_260_p2;
reg   [42:0] r_V_190_reg_2331;
wire   [53:0] r_V_191_fu_263_p2;
reg   [53:0] r_V_191_reg_2335;
wire   [42:0] r_V_192_fu_250_p2;
reg   [42:0] r_V_192_reg_2339;
wire   [42:0] r_V_193_fu_244_p2;
reg   [42:0] r_V_193_reg_2343;
wire   [53:0] r_V_194_fu_243_p2;
reg   [53:0] r_V_194_reg_2347;
wire   [53:0] r_V_195_fu_248_p2;
reg   [53:0] r_V_195_reg_2351;
wire   [42:0] r_V_fu_247_p2;
reg   [42:0] r_V_reg_2675;
wire   [41:0] r_V_196_fu_258_p2;
reg   [41:0] r_V_196_reg_2679;
wire   [43:0] r_V_197_fu_245_p2;
reg   [43:0] r_V_197_reg_2683;
wire   [44:0] r_V_198_fu_265_p2;
reg   [44:0] r_V_198_reg_2687;
wire   [53:0] r_V_199_fu_255_p2;
reg   [53:0] r_V_199_reg_2691;
wire   [40:0] r_V_201_fu_257_p2;
reg   [40:0] r_V_201_reg_2695;
wire   [53:0] r_V_202_fu_252_p2;
reg   [53:0] r_V_202_reg_2699;
wire   [53:0] r_V_203_fu_253_p2;
reg   [53:0] r_V_203_reg_2703;
reg   [0:0] p_Result_s_reg_10769;
reg   [0:0] p_Result_807_reg_10775;
wire  signed [19:0] p_Val2_807_fu_2783_p2;
reg  signed [19:0] p_Val2_807_reg_10781;
reg   [0:0] p_Result_808_reg_10786;
reg   [0:0] Range2_all_ones_reg_10793;
reg   [0:0] p_Result_809_reg_10800;
reg   [0:0] p_Result_810_reg_10806;
wire  signed [20:0] p_Val2_810_fu_2847_p2;
reg  signed [20:0] p_Val2_810_reg_10812;
reg   [0:0] p_Result_811_reg_10817;
reg   [0:0] Range2_all_ones_159_reg_10824;
reg   [0:0] p_Result_812_reg_10831;
reg   [0:0] p_Result_813_reg_10837;
wire   [31:0] p_Val2_813_fu_2907_p2;
reg   [31:0] p_Val2_813_reg_10843;
reg   [0:0] p_Result_814_reg_10848;
reg   [0:0] Range2_all_ones_160_reg_10855;
reg   [0:0] p_Result_815_reg_10862;
reg   [0:0] p_Result_816_reg_10868;
wire  signed [20:0] p_Val2_816_fu_2971_p2;
reg  signed [20:0] p_Val2_816_reg_10874;
reg   [0:0] p_Result_817_reg_10879;
reg   [0:0] Range2_all_ones_161_reg_10886;
reg   [0:0] p_Result_818_reg_10893;
reg   [0:0] p_Result_819_reg_10899;
wire  signed [23:0] p_Val2_819_fu_3035_p2;
reg  signed [23:0] p_Val2_819_reg_10905;
reg   [0:0] p_Result_820_reg_10910;
reg   [0:0] Range2_all_ones_162_reg_10917;
reg   [0:0] p_Result_821_reg_10924;
reg   [0:0] p_Result_822_reg_10930;
wire  signed [19:0] p_Val2_822_fu_3099_p2;
reg  signed [19:0] p_Val2_822_reg_10936;
reg   [0:0] p_Result_823_reg_10941;
reg   [0:0] Range2_all_ones_163_reg_10948;
reg   [0:0] p_Result_824_reg_10955;
reg   [0:0] p_Result_825_reg_10961;
wire  signed [19:0] p_Val2_825_fu_3163_p2;
reg  signed [19:0] p_Val2_825_reg_10967;
reg   [0:0] p_Result_826_reg_10972;
reg   [0:0] Range2_all_ones_164_reg_10979;
reg   [0:0] p_Result_827_reg_10986;
reg   [0:0] p_Result_828_reg_10992;
wire  signed [30:0] p_Val2_828_fu_3227_p2;
reg  signed [30:0] p_Val2_828_reg_10998;
reg   [0:0] p_Result_829_reg_11003;
reg   [0:0] Range2_all_ones_165_reg_11010;
reg   [0:0] p_Result_830_reg_11017;
reg   [0:0] p_Result_831_reg_11023;
wire  signed [30:0] p_Val2_831_fu_3291_p2;
reg  signed [30:0] p_Val2_831_reg_11029;
reg   [0:0] p_Result_832_reg_11034;
reg   [0:0] Range2_all_ones_166_reg_11041;
reg   [0:0] p_Result_833_reg_11048;
reg   [16:0] p_Val2_833_reg_11054;
reg   [0:0] p_Result_834_reg_11059;
reg   [0:0] tmp_1338_reg_11065;
reg   [0:0] Range2_all_ones_167_reg_11070;
reg   [0:0] p_Result_836_reg_11077;
reg   [18:0] p_Val2_836_reg_11083;
reg   [0:0] p_Result_837_reg_11088;
reg   [0:0] tmp_1344_reg_11094;
reg   [0:0] Range2_all_ones_168_reg_11099;
reg   [0:0] p_Result_839_reg_11106;
reg   [20:0] p_Val2_839_reg_11112;
reg   [0:0] p_Result_840_reg_11117;
reg   [0:0] tmp_1350_reg_11123;
reg   [0:0] Range2_all_ones_169_reg_11128;
reg   [0:0] p_Result_842_reg_11135;
reg   [18:0] p_Val2_842_reg_11141;
reg   [0:0] p_Result_843_reg_11146;
reg   [0:0] tmp_1356_reg_11152;
reg   [0:0] Range2_all_ones_170_reg_11157;
reg   [0:0] p_Result_845_reg_11164;
reg   [29:0] p_Val2_845_reg_11170;
reg   [0:0] p_Result_846_reg_11175;
reg   [0:0] tmp_1362_reg_11181;
reg   [0:0] Range2_all_ones_171_reg_11186;
reg   [0:0] p_Result_848_reg_11193;
reg   [18:0] p_Val2_848_reg_11199;
reg   [0:0] p_Result_849_reg_11204;
reg   [0:0] tmp_1368_reg_11210;
reg   [0:0] Range2_all_ones_172_reg_11215;
reg   [0:0] p_Result_851_reg_11222;
reg   [18:0] p_Val2_851_reg_11228;
reg   [0:0] p_Result_852_reg_11233;
reg   [0:0] tmp_1374_reg_11239;
reg   [0:0] Range2_all_ones_173_reg_11244;
reg   [0:0] p_Result_854_reg_11251;
reg   [29:0] p_Val2_854_reg_11257;
reg   [0:0] p_Result_855_reg_11262;
reg   [0:0] tmp_1380_reg_11268;
reg   [0:0] Range2_all_ones_174_reg_11273;
reg   [0:0] p_Result_857_reg_11280;
reg   [29:0] p_Val2_857_reg_11286;
reg   [0:0] p_Result_858_reg_11291;
reg   [0:0] tmp_1386_reg_11297;
reg   [0:0] Range2_all_ones_175_reg_11302;
wire  signed [31:0] a_V_2_fu_3726_p4;
reg  signed [31:0] a_V_2_reg_11309;
wire  signed [15:0] p_Val2_876_fu_3844_p2;
reg  signed [15:0] p_Val2_876_reg_11319;
reg  signed [15:0] p_Val2_876_reg_11319_pp0_iter1_reg;
wire   [0:0] overflow_345_fu_3946_p2;
reg   [0:0] overflow_345_reg_11324;
reg   [0:0] overflow_345_reg_11324_pp0_iter1_reg;
wire   [0:0] or_ln346_183_fu_3976_p2;
reg   [0:0] or_ln346_183_reg_11329;
reg   [0:0] or_ln346_183_reg_11329_pp0_iter1_reg;
reg   [0:0] p_Result_860_reg_11334;
reg   [18:0] p_Val2_860_reg_11340;
reg   [0:0] p_Result_861_reg_11345;
reg   [0:0] tmp_1392_reg_11351;
reg   [0:0] Range2_all_ones_176_reg_11356;
reg   [0:0] p_Result_863_reg_11363;
reg   [17:0] p_Val2_863_reg_11369;
reg   [0:0] p_Result_864_reg_11374;
reg   [0:0] tmp_1398_reg_11380;
reg   [0:0] Range2_all_ones_177_reg_11385;
reg   [0:0] p_Result_866_reg_11392;
reg   [19:0] p_Val2_866_reg_11398;
reg   [0:0] p_Result_867_reg_11403;
reg   [0:0] tmp_1404_reg_11409;
reg   [0:0] Range2_all_ones_178_reg_11414;
reg   [0:0] p_Result_869_reg_11421;
reg   [20:0] p_Val2_869_reg_11427;
reg   [0:0] p_Result_870_reg_11432;
reg   [0:0] tmp_1410_reg_11438;
reg   [0:0] Range2_all_ones_179_reg_11443;
reg   [0:0] p_Result_872_reg_11450;
reg   [29:0] p_Val2_872_reg_11456;
reg   [0:0] p_Result_873_reg_11461;
reg   [0:0] tmp_1416_reg_11467;
reg   [0:0] Range2_all_ones_180_reg_11472;
reg   [0:0] p_Result_878_reg_11479;
reg   [16:0] p_Val2_878_reg_11485;
reg   [0:0] p_Result_879_reg_11490;
reg   [0:0] tmp_1428_reg_11496;
reg   [0:0] Range2_all_ones_182_reg_11501;
reg   [0:0] p_Result_881_reg_11508;
reg   [29:0] p_Val2_881_reg_11514;
reg   [0:0] p_Result_882_reg_11519;
reg   [0:0] tmp_1434_reg_11525;
reg   [0:0] Range2_all_ones_183_reg_11530;
reg   [0:0] p_Result_884_reg_11537;
reg   [29:0] p_Val2_884_reg_11543;
reg   [0:0] p_Result_885_reg_11548;
reg   [0:0] tmp_1440_reg_11554;
reg   [0:0] Range2_all_ones_184_reg_11559;
wire  signed [31:0] lhs_151_fu_7782_p3;
reg  signed [31:0] lhs_151_reg_11566;
wire  signed [31:0] lhs_152_fu_7884_p3;
reg  signed [31:0] lhs_152_reg_11572;
wire  signed [31:0] lhs_153_fu_7986_p3;
reg  signed [31:0] lhs_153_reg_11578;
wire  signed [31:0] lhs_154_fu_8088_p3;
reg  signed [31:0] lhs_154_reg_11584;
wire  signed [31:0] lhs_155_fu_8190_p3;
reg  signed [31:0] lhs_155_reg_11590;
wire  signed [31:0] lhs_156_fu_8292_p3;
reg  signed [31:0] lhs_156_reg_11596;
wire  signed [31:0] lhs_157_fu_8394_p3;
reg  signed [31:0] lhs_157_reg_11602;
wire  signed [31:0] lhs_158_fu_8496_p3;
reg  signed [31:0] lhs_158_reg_11608;
wire  signed [31:0] lhs_159_fu_8598_p3;
reg  signed [31:0] lhs_159_reg_11614;
wire  signed [31:0] r_V_183_fu_240_p0;
wire  signed [42:0] sext_ln70_93_fu_2734_p1;
wire   [10:0] r_V_183_fu_240_p1;
wire    ap_block_pp0_stage0;
wire  signed [12:0] r_V_189_fu_242_p1;
wire  signed [31:0] r_V_194_fu_243_p0;
wire  signed [53:0] sext_ln70_94_fu_3323_p1;
wire  signed [22:0] r_V_194_fu_243_p1;
wire  signed [31:0] r_V_193_fu_244_p0;
wire  signed [42:0] sext_ln70_96_fu_3335_p1;
wire  signed [10:0] r_V_193_fu_244_p1;
wire   [11:0] r_V_197_fu_245_p1;
wire  signed [31:0] r_V_186_fu_246_p0;
wire  signed [53:0] sext_ln70_fu_2712_p1;
wire   [22:0] r_V_186_fu_246_p1;
wire  signed [10:0] r_V_fu_247_p1;
wire  signed [31:0] r_V_195_fu_248_p0;
wire  signed [22:0] r_V_195_fu_248_p1;
wire  signed [31:0] r_V_184_fu_249_p0;
wire   [10:0] r_V_184_fu_249_p1;
wire  signed [31:0] r_V_192_fu_250_p0;
wire   [10:0] r_V_192_fu_250_p1;
wire   [25:0] r_V_180_fu_251_p1;
wire  signed [31:0] r_V_202_fu_252_p0;
wire  signed [53:0] sext_ln70_100_fu_6448_p1;
wire   [22:0] r_V_202_fu_252_p1;
wire  signed [31:0] r_V_203_fu_253_p0;
wire   [22:0] r_V_203_fu_253_p1;
wire  signed [31:0] r_V_178_fu_254_p0;
wire  signed [10:0] r_V_178_fu_254_p1;
wire  signed [31:0] r_V_199_fu_255_p0;
wire  signed [22:0] r_V_199_fu_255_p1;
wire  signed [31:0] r_V_181_fu_256_p0;
wire  signed [43:0] sext_ln70_92_fu_2728_p1;
wire  signed [11:0] r_V_181_fu_256_p1;
wire  signed [8:0] r_V_201_fu_257_p1;
wire  signed [9:0] r_V_196_fu_258_p1;
wire  signed [31:0] r_V_185_fu_259_p0;
wire   [22:0] r_V_185_fu_259_p1;
wire  signed [31:0] r_V_190_fu_260_p0;
wire   [10:0] r_V_190_fu_260_p1;
wire  signed [31:0] r_V_188_fu_261_p0;
wire   [10:0] r_V_188_fu_261_p1;
wire  signed [31:0] r_V_179_fu_262_p0;
wire  signed [11:0] r_V_179_fu_262_p1;
wire  signed [31:0] r_V_191_fu_263_p0;
wire   [22:0] r_V_191_fu_263_p1;
wire   [14:0] r_V_182_fu_264_p1;
wire  signed [12:0] r_V_198_fu_265_p1;
wire  signed [8:0] r_V_187_fu_266_p1;
wire  signed [31:0] a_V_fu_2708_p1;
wire   [18:0] p_Val2_806_fu_2749_p4;
wire   [0:0] tmp_fu_2771_p3;
wire   [19:0] zext_ln377_fu_2779_p1;
wire  signed [19:0] sext_ln823_fu_2759_p1;
wire   [19:0] p_Val2_809_fu_2813_p4;
wire   [0:0] tmp_1290_fu_2835_p3;
wire   [20:0] zext_ln377_161_fu_2843_p1;
wire  signed [20:0] sext_ln823_153_fu_2823_p1;
wire   [0:0] tmp_1296_fu_2895_p3;
wire   [31:0] zext_ln377_162_fu_2903_p1;
wire   [31:0] p_Val2_812_fu_2877_p4;
wire   [19:0] p_Val2_815_fu_2937_p4;
wire   [0:0] tmp_1302_fu_2959_p3;
wire   [20:0] zext_ln377_163_fu_2967_p1;
wire  signed [20:0] sext_ln823_154_fu_2947_p1;
wire   [22:0] p_Val2_818_fu_3001_p4;
wire   [0:0] tmp_1308_fu_3023_p3;
wire   [23:0] zext_ln377_164_fu_3031_p1;
wire  signed [23:0] sext_ln823_155_fu_3011_p1;
wire   [18:0] p_Val2_821_fu_3065_p4;
wire   [0:0] tmp_1314_fu_3087_p3;
wire   [19:0] zext_ln377_165_fu_3095_p1;
wire  signed [19:0] sext_ln823_156_fu_3075_p1;
wire   [18:0] p_Val2_824_fu_3129_p4;
wire   [0:0] tmp_1320_fu_3151_p3;
wire   [19:0] zext_ln377_166_fu_3159_p1;
wire  signed [19:0] sext_ln823_157_fu_3139_p1;
wire   [29:0] p_Val2_827_fu_3193_p4;
wire   [0:0] tmp_1326_fu_3215_p3;
wire   [30:0] zext_ln377_167_fu_3223_p1;
wire  signed [30:0] sext_ln823_158_fu_3203_p1;
wire   [29:0] p_Val2_830_fu_3257_p4;
wire   [0:0] tmp_1332_fu_3279_p3;
wire   [30:0] zext_ln377_168_fu_3287_p1;
wire  signed [30:0] sext_ln823_159_fu_3267_p1;
wire  signed [31:0] a_V_1_fu_3313_p4;
wire   [31:0] tmp288_fu_3750_p4;
wire   [37:0] shl_ln_fu_3760_p3;
wire   [17:0] tmp_s_fu_3772_p4;
wire  signed [38:0] sext_ln1273_fu_3768_p1;
wire  signed [38:0] sext_ln70_99_fu_3746_p1;
wire   [38:0] r_V_200_fu_3790_p2;
wire   [14:0] p_Val2_875_fu_3804_p4;
wire   [23:0] trunc_ln7_fu_3782_p3;
wire   [23:0] a_V_2_cast_fu_3736_p4;
wire   [23:0] add_ln823_fu_3818_p2;
wire   [0:0] tmp_1422_fu_3832_p3;
wire   [15:0] zext_ln377_183_fu_3840_p1;
wire  signed [15:0] sext_ln823_174_fu_3814_p1;
wire   [0:0] p_Result_877_fu_3850_p3;
wire   [0:0] p_Result_876_fu_3824_p3;
wire   [0:0] xor_ln896_530_fu_3858_p2;
wire   [0:0] xor_ln888_365_fu_3878_p2;
wire   [0:0] Range2_all_ones_181_fu_3870_p3;
wire   [0:0] or_ln888_183_fu_3884_p2;
wire   [0:0] tmp_1425_fu_3896_p3;
wire   [0:0] xor_ln890_181_fu_3904_p2;
wire   [0:0] or_ln890_183_fu_3910_p2;
wire   [0:0] carry_366_fu_3864_p2;
wire   [0:0] deleted_zeros_180_fu_3890_p2;
wire   [0:0] xor_ln895_530_fu_3928_p2;
wire   [0:0] p_Result_875_fu_3796_p3;
wire   [0:0] or_ln895_183_fu_3934_p2;
wire   [0:0] xor_ln895_531_fu_3940_p2;
wire   [0:0] deleted_ones_345_fu_3916_p2;
wire   [0:0] xor_ln896_531_fu_3952_p2;
wire   [0:0] and_ln891_183_fu_3922_p2;
wire   [0:0] or_ln896_183_fu_3958_p2;
wire   [0:0] xor_ln896_589_fu_3964_p2;
wire   [0:0] underflow_345_fu_3970_p2;
wire   [0:0] xor_ln896_fu_3985_p2;
wire   [0:0] xor_ln888_fu_3995_p2;
wire   [0:0] or_ln888_fu_4000_p2;
wire   [0:0] tmp_1287_fu_4010_p3;
wire   [0:0] xor_ln890_fu_4018_p2;
wire   [0:0] or_ln890_fu_4024_p2;
wire   [0:0] carry_320_fu_3990_p2;
wire   [0:0] deleted_zeros_fu_4005_p2;
wire   [0:0] xor_ln895_fu_4040_p2;
wire   [0:0] or_ln895_fu_4046_p2;
wire   [0:0] xor_ln895_485_fu_4051_p2;
wire   [0:0] deleted_ones_fu_4030_p2;
wire   [0:0] xor_ln896_485_fu_4062_p2;
wire   [0:0] and_ln891_fu_4035_p2;
wire   [0:0] or_ln896_fu_4068_p2;
wire   [0:0] xor_ln896_566_fu_4074_p2;
wire   [0:0] overflow_fu_4056_p2;
wire   [0:0] underflow_fu_4080_p2;
wire   [0:0] or_ln346_fu_4093_p2;
wire   [31:0] select_ln346_243_fu_4085_p3;
wire  signed [31:0] sext_ln856_fu_3982_p1;
wire   [0:0] xor_ln896_486_fu_4110_p2;
wire   [0:0] xor_ln888_321_fu_4120_p2;
wire   [0:0] or_ln888_161_fu_4125_p2;
wire   [0:0] tmp_1293_fu_4135_p3;
wire   [0:0] xor_ln890_159_fu_4143_p2;
wire   [0:0] or_ln890_161_fu_4149_p2;
wire   [0:0] carry_322_fu_4115_p2;
wire   [0:0] deleted_zeros_158_fu_4130_p2;
wire   [0:0] xor_ln895_486_fu_4165_p2;
wire   [0:0] or_ln895_161_fu_4171_p2;
wire   [0:0] xor_ln895_487_fu_4176_p2;
wire   [0:0] deleted_ones_323_fu_4155_p2;
wire   [0:0] xor_ln896_487_fu_4187_p2;
wire   [0:0] and_ln891_161_fu_4160_p2;
wire   [0:0] or_ln896_161_fu_4193_p2;
wire   [0:0] xor_ln896_567_fu_4199_p2;
wire   [0:0] overflow_323_fu_4181_p2;
wire   [0:0] underflow_323_fu_4205_p2;
wire   [0:0] or_ln346_161_fu_4218_p2;
wire   [31:0] select_ln346_244_fu_4210_p3;
wire  signed [31:0] sext_ln856_153_fu_4107_p1;
wire   [0:0] xor_ln896_488_fu_4232_p2;
wire   [0:0] xor_ln888_323_fu_4242_p2;
wire   [0:0] or_ln888_162_fu_4247_p2;
wire   [0:0] tmp_1299_fu_4257_p3;
wire   [0:0] xor_ln890_160_fu_4265_p2;
wire   [0:0] or_ln890_162_fu_4271_p2;
wire   [0:0] carry_324_fu_4237_p2;
wire   [0:0] deleted_zeros_159_fu_4252_p2;
wire   [0:0] xor_ln895_488_fu_4287_p2;
wire   [0:0] or_ln895_162_fu_4293_p2;
wire   [0:0] xor_ln895_489_fu_4298_p2;
wire   [0:0] deleted_ones_324_fu_4277_p2;
wire   [0:0] xor_ln896_489_fu_4309_p2;
wire   [0:0] and_ln891_162_fu_4282_p2;
wire   [0:0] or_ln896_162_fu_4315_p2;
wire   [0:0] xor_ln896_568_fu_4321_p2;
wire   [0:0] overflow_324_fu_4303_p2;
wire   [0:0] underflow_324_fu_4327_p2;
wire   [0:0] or_ln346_162_fu_4340_p2;
wire   [31:0] select_ln346_245_fu_4332_p3;
wire   [0:0] xor_ln896_490_fu_4356_p2;
wire   [0:0] xor_ln888_325_fu_4366_p2;
wire   [0:0] or_ln888_163_fu_4371_p2;
wire   [0:0] tmp_1305_fu_4381_p3;
wire   [0:0] xor_ln890_161_fu_4389_p2;
wire   [0:0] or_ln890_163_fu_4395_p2;
wire   [0:0] carry_326_fu_4361_p2;
wire   [0:0] deleted_zeros_160_fu_4376_p2;
wire   [0:0] xor_ln895_490_fu_4411_p2;
wire   [0:0] or_ln895_163_fu_4417_p2;
wire   [0:0] xor_ln895_491_fu_4422_p2;
wire   [0:0] deleted_ones_325_fu_4401_p2;
wire   [0:0] xor_ln896_491_fu_4433_p2;
wire   [0:0] and_ln891_163_fu_4406_p2;
wire   [0:0] or_ln896_163_fu_4439_p2;
wire   [0:0] xor_ln896_569_fu_4445_p2;
wire   [0:0] overflow_325_fu_4427_p2;
wire   [0:0] underflow_325_fu_4451_p2;
wire   [0:0] or_ln346_163_fu_4464_p2;
wire   [31:0] select_ln346_246_fu_4456_p3;
wire  signed [31:0] sext_ln856_154_fu_4353_p1;
wire   [0:0] xor_ln896_492_fu_4481_p2;
wire   [0:0] xor_ln888_327_fu_4491_p2;
wire   [0:0] or_ln888_164_fu_4496_p2;
wire   [0:0] tmp_1311_fu_4506_p3;
wire   [0:0] xor_ln890_162_fu_4514_p2;
wire   [0:0] or_ln890_164_fu_4520_p2;
wire   [0:0] carry_328_fu_4486_p2;
wire   [0:0] deleted_zeros_161_fu_4501_p2;
wire   [0:0] xor_ln895_492_fu_4536_p2;
wire   [0:0] or_ln895_164_fu_4542_p2;
wire   [0:0] xor_ln895_493_fu_4547_p2;
wire   [0:0] deleted_ones_326_fu_4526_p2;
wire   [0:0] xor_ln896_493_fu_4558_p2;
wire   [0:0] and_ln891_164_fu_4531_p2;
wire   [0:0] or_ln896_164_fu_4564_p2;
wire   [0:0] xor_ln896_570_fu_4570_p2;
wire   [0:0] overflow_326_fu_4552_p2;
wire   [0:0] underflow_326_fu_4576_p2;
wire   [0:0] or_ln346_164_fu_4589_p2;
wire   [31:0] select_ln346_247_fu_4581_p3;
wire  signed [31:0] sext_ln856_155_fu_4478_p1;
wire   [0:0] xor_ln896_494_fu_4606_p2;
wire   [0:0] xor_ln888_329_fu_4616_p2;
wire   [0:0] or_ln888_165_fu_4621_p2;
wire   [0:0] tmp_1317_fu_4631_p3;
wire   [0:0] xor_ln890_163_fu_4639_p2;
wire   [0:0] or_ln890_165_fu_4645_p2;
wire   [0:0] carry_330_fu_4611_p2;
wire   [0:0] deleted_zeros_162_fu_4626_p2;
wire   [0:0] xor_ln895_494_fu_4661_p2;
wire   [0:0] or_ln895_165_fu_4667_p2;
wire   [0:0] xor_ln895_495_fu_4672_p2;
wire   [0:0] deleted_ones_327_fu_4651_p2;
wire   [0:0] xor_ln896_495_fu_4683_p2;
wire   [0:0] and_ln891_165_fu_4656_p2;
wire   [0:0] or_ln896_165_fu_4689_p2;
wire   [0:0] xor_ln896_571_fu_4695_p2;
wire   [0:0] overflow_327_fu_4677_p2;
wire   [0:0] underflow_327_fu_4701_p2;
wire   [0:0] or_ln346_165_fu_4714_p2;
wire   [31:0] select_ln346_248_fu_4706_p3;
wire  signed [31:0] sext_ln856_156_fu_4603_p1;
wire   [0:0] xor_ln896_496_fu_4731_p2;
wire   [0:0] xor_ln888_331_fu_4741_p2;
wire   [0:0] or_ln888_166_fu_4746_p2;
wire   [0:0] tmp_1323_fu_4756_p3;
wire   [0:0] xor_ln890_164_fu_4764_p2;
wire   [0:0] or_ln890_166_fu_4770_p2;
wire   [0:0] carry_332_fu_4736_p2;
wire   [0:0] deleted_zeros_163_fu_4751_p2;
wire   [0:0] xor_ln895_496_fu_4786_p2;
wire   [0:0] or_ln895_166_fu_4792_p2;
wire   [0:0] xor_ln895_497_fu_4797_p2;
wire   [0:0] deleted_ones_328_fu_4776_p2;
wire   [0:0] xor_ln896_497_fu_4808_p2;
wire   [0:0] and_ln891_166_fu_4781_p2;
wire   [0:0] or_ln896_166_fu_4814_p2;
wire   [0:0] xor_ln896_572_fu_4820_p2;
wire   [0:0] overflow_328_fu_4802_p2;
wire   [0:0] underflow_328_fu_4826_p2;
wire   [0:0] or_ln346_166_fu_4839_p2;
wire   [31:0] select_ln346_249_fu_4831_p3;
wire  signed [31:0] sext_ln856_157_fu_4728_p1;
wire   [0:0] xor_ln896_498_fu_4856_p2;
wire   [0:0] xor_ln888_333_fu_4866_p2;
wire   [0:0] or_ln888_167_fu_4871_p2;
wire   [0:0] tmp_1329_fu_4881_p3;
wire   [0:0] xor_ln890_165_fu_4889_p2;
wire   [0:0] or_ln890_167_fu_4895_p2;
wire   [0:0] carry_334_fu_4861_p2;
wire   [0:0] deleted_zeros_164_fu_4876_p2;
wire   [0:0] xor_ln895_498_fu_4911_p2;
wire   [0:0] or_ln895_167_fu_4917_p2;
wire   [0:0] xor_ln895_499_fu_4922_p2;
wire   [0:0] deleted_ones_329_fu_4901_p2;
wire   [0:0] xor_ln896_499_fu_4933_p2;
wire   [0:0] and_ln891_167_fu_4906_p2;
wire   [0:0] or_ln896_167_fu_4939_p2;
wire   [0:0] xor_ln896_573_fu_4945_p2;
wire   [0:0] overflow_329_fu_4927_p2;
wire   [0:0] underflow_329_fu_4951_p2;
wire   [0:0] or_ln346_167_fu_4964_p2;
wire   [31:0] select_ln346_250_fu_4956_p3;
wire  signed [31:0] sext_ln856_158_fu_4853_p1;
wire   [0:0] xor_ln896_500_fu_4981_p2;
wire   [0:0] xor_ln888_335_fu_4991_p2;
wire   [0:0] or_ln888_168_fu_4996_p2;
wire   [0:0] tmp_1335_fu_5006_p3;
wire   [0:0] xor_ln890_166_fu_5014_p2;
wire   [0:0] or_ln890_168_fu_5020_p2;
wire   [0:0] carry_336_fu_4986_p2;
wire   [0:0] deleted_zeros_165_fu_5001_p2;
wire   [0:0] xor_ln895_500_fu_5036_p2;
wire   [0:0] or_ln895_168_fu_5042_p2;
wire   [0:0] xor_ln895_501_fu_5047_p2;
wire   [0:0] deleted_ones_330_fu_5026_p2;
wire   [0:0] xor_ln896_501_fu_5058_p2;
wire   [0:0] and_ln891_168_fu_5031_p2;
wire   [0:0] or_ln896_168_fu_5064_p2;
wire   [0:0] xor_ln896_574_fu_5070_p2;
wire   [0:0] overflow_330_fu_5052_p2;
wire   [0:0] underflow_330_fu_5076_p2;
wire   [0:0] or_ln346_168_fu_5089_p2;
wire   [31:0] select_ln346_251_fu_5081_p3;
wire  signed [31:0] sext_ln856_159_fu_4978_p1;
wire   [17:0] zext_ln377_169_fu_5106_p1;
wire  signed [17:0] sext_ln823_160_fu_5103_p1;
wire  signed [17:0] p_Val2_834_fu_5109_p2;
wire   [0:0] p_Result_835_fu_5119_p3;
wire   [0:0] xor_ln896_502_fu_5127_p2;
wire   [0:0] xor_ln888_337_fu_5138_p2;
wire   [0:0] or_ln888_169_fu_5143_p2;
wire   [0:0] tmp_1341_fu_5154_p3;
wire   [0:0] xor_ln890_167_fu_5162_p2;
wire   [0:0] or_ln890_169_fu_5168_p2;
wire   [0:0] carry_338_fu_5133_p2;
wire   [0:0] deleted_zeros_166_fu_5149_p2;
wire   [0:0] xor_ln895_502_fu_5184_p2;
wire   [0:0] or_ln895_169_fu_5190_p2;
wire   [0:0] xor_ln895_503_fu_5196_p2;
wire   [0:0] deleted_ones_331_fu_5174_p2;
wire   [0:0] xor_ln896_503_fu_5207_p2;
wire   [0:0] and_ln891_169_fu_5179_p2;
wire   [0:0] or_ln896_169_fu_5213_p2;
wire   [0:0] xor_ln896_575_fu_5219_p2;
wire   [0:0] overflow_331_fu_5201_p2;
wire   [0:0] underflow_331_fu_5225_p2;
wire   [0:0] or_ln346_169_fu_5238_p2;
wire   [31:0] select_ln346_252_fu_5230_p3;
wire  signed [31:0] sext_ln856_160_fu_5115_p1;
wire   [19:0] zext_ln377_170_fu_5255_p1;
wire  signed [19:0] sext_ln823_161_fu_5252_p1;
wire  signed [19:0] p_Val2_837_fu_5258_p2;
wire   [0:0] p_Result_838_fu_5268_p3;
wire   [0:0] xor_ln896_504_fu_5276_p2;
wire   [0:0] xor_ln888_339_fu_5287_p2;
wire   [0:0] or_ln888_170_fu_5292_p2;
wire   [0:0] tmp_1347_fu_5303_p3;
wire   [0:0] xor_ln890_168_fu_5311_p2;
wire   [0:0] or_ln890_170_fu_5317_p2;
wire   [0:0] carry_340_fu_5282_p2;
wire   [0:0] deleted_zeros_167_fu_5298_p2;
wire   [0:0] xor_ln895_504_fu_5333_p2;
wire   [0:0] or_ln895_170_fu_5339_p2;
wire   [0:0] xor_ln895_505_fu_5345_p2;
wire   [0:0] deleted_ones_332_fu_5323_p2;
wire   [0:0] xor_ln896_505_fu_5356_p2;
wire   [0:0] and_ln891_170_fu_5328_p2;
wire   [0:0] or_ln896_170_fu_5362_p2;
wire   [0:0] xor_ln896_576_fu_5368_p2;
wire   [0:0] overflow_332_fu_5350_p2;
wire   [0:0] underflow_332_fu_5374_p2;
wire   [0:0] or_ln346_170_fu_5387_p2;
wire   [31:0] select_ln346_253_fu_5379_p3;
wire  signed [31:0] sext_ln856_161_fu_5264_p1;
wire   [21:0] zext_ln377_171_fu_5404_p1;
wire  signed [21:0] sext_ln823_162_fu_5401_p1;
wire  signed [21:0] p_Val2_840_fu_5407_p2;
wire   [0:0] p_Result_841_fu_5417_p3;
wire   [0:0] xor_ln896_506_fu_5425_p2;
wire   [0:0] xor_ln888_341_fu_5436_p2;
wire   [0:0] or_ln888_171_fu_5441_p2;
wire   [0:0] tmp_1353_fu_5452_p3;
wire   [0:0] xor_ln890_169_fu_5460_p2;
wire   [0:0] or_ln890_171_fu_5466_p2;
wire   [0:0] carry_342_fu_5431_p2;
wire   [0:0] deleted_zeros_168_fu_5447_p2;
wire   [0:0] xor_ln895_506_fu_5482_p2;
wire   [0:0] or_ln895_171_fu_5488_p2;
wire   [0:0] xor_ln895_507_fu_5494_p2;
wire   [0:0] deleted_ones_333_fu_5472_p2;
wire   [0:0] xor_ln896_507_fu_5505_p2;
wire   [0:0] and_ln891_171_fu_5477_p2;
wire   [0:0] or_ln896_171_fu_5511_p2;
wire   [0:0] xor_ln896_577_fu_5517_p2;
wire   [0:0] overflow_333_fu_5499_p2;
wire   [0:0] underflow_333_fu_5523_p2;
wire   [0:0] or_ln346_171_fu_5536_p2;
wire   [31:0] select_ln346_254_fu_5528_p3;
wire  signed [31:0] sext_ln856_162_fu_5413_p1;
wire   [19:0] zext_ln377_172_fu_5553_p1;
wire  signed [19:0] sext_ln823_163_fu_5550_p1;
wire  signed [19:0] p_Val2_843_fu_5556_p2;
wire   [0:0] p_Result_844_fu_5566_p3;
wire   [0:0] xor_ln896_508_fu_5574_p2;
wire   [0:0] xor_ln888_343_fu_5585_p2;
wire   [0:0] or_ln888_172_fu_5590_p2;
wire   [0:0] tmp_1359_fu_5601_p3;
wire   [0:0] xor_ln890_170_fu_5609_p2;
wire   [0:0] or_ln890_172_fu_5615_p2;
wire   [0:0] carry_344_fu_5580_p2;
wire   [0:0] deleted_zeros_169_fu_5596_p2;
wire   [0:0] xor_ln895_508_fu_5631_p2;
wire   [0:0] or_ln895_172_fu_5637_p2;
wire   [0:0] xor_ln895_509_fu_5643_p2;
wire   [0:0] deleted_ones_334_fu_5621_p2;
wire   [0:0] xor_ln896_509_fu_5654_p2;
wire   [0:0] and_ln891_172_fu_5626_p2;
wire   [0:0] or_ln896_172_fu_5660_p2;
wire   [0:0] xor_ln896_578_fu_5666_p2;
wire   [0:0] overflow_334_fu_5648_p2;
wire   [0:0] underflow_334_fu_5672_p2;
wire   [0:0] or_ln346_172_fu_5685_p2;
wire   [31:0] select_ln346_255_fu_5677_p3;
wire  signed [31:0] sext_ln856_163_fu_5562_p1;
wire   [30:0] zext_ln377_173_fu_5702_p1;
wire  signed [30:0] sext_ln823_164_fu_5699_p1;
wire  signed [30:0] p_Val2_846_fu_5705_p2;
wire   [0:0] p_Result_847_fu_5715_p3;
wire   [0:0] xor_ln896_510_fu_5723_p2;
wire   [0:0] xor_ln888_345_fu_5734_p2;
wire   [0:0] or_ln888_173_fu_5739_p2;
wire   [0:0] tmp_1365_fu_5750_p3;
wire   [0:0] xor_ln890_171_fu_5758_p2;
wire   [0:0] or_ln890_173_fu_5764_p2;
wire   [0:0] carry_346_fu_5729_p2;
wire   [0:0] deleted_zeros_170_fu_5745_p2;
wire   [0:0] xor_ln895_510_fu_5780_p2;
wire   [0:0] or_ln895_173_fu_5786_p2;
wire   [0:0] xor_ln895_511_fu_5792_p2;
wire   [0:0] deleted_ones_335_fu_5770_p2;
wire   [0:0] xor_ln896_511_fu_5803_p2;
wire   [0:0] and_ln891_173_fu_5775_p2;
wire   [0:0] or_ln896_173_fu_5809_p2;
wire   [0:0] xor_ln896_579_fu_5815_p2;
wire   [0:0] overflow_335_fu_5797_p2;
wire   [0:0] underflow_335_fu_5821_p2;
wire   [0:0] or_ln346_173_fu_5834_p2;
wire   [31:0] select_ln346_256_fu_5826_p3;
wire  signed [31:0] sext_ln856_164_fu_5711_p1;
wire   [19:0] zext_ln377_174_fu_5851_p1;
wire  signed [19:0] sext_ln823_165_fu_5848_p1;
wire  signed [19:0] p_Val2_849_fu_5854_p2;
wire   [0:0] p_Result_850_fu_5864_p3;
wire   [0:0] xor_ln896_512_fu_5872_p2;
wire   [0:0] xor_ln888_347_fu_5883_p2;
wire   [0:0] or_ln888_174_fu_5888_p2;
wire   [0:0] tmp_1371_fu_5899_p3;
wire   [0:0] xor_ln890_172_fu_5907_p2;
wire   [0:0] or_ln890_174_fu_5913_p2;
wire   [0:0] carry_348_fu_5878_p2;
wire   [0:0] deleted_zeros_171_fu_5894_p2;
wire   [0:0] xor_ln895_512_fu_5929_p2;
wire   [0:0] or_ln895_174_fu_5935_p2;
wire   [0:0] xor_ln895_513_fu_5941_p2;
wire   [0:0] deleted_ones_336_fu_5919_p2;
wire   [0:0] xor_ln896_513_fu_5952_p2;
wire   [0:0] and_ln891_174_fu_5924_p2;
wire   [0:0] or_ln896_174_fu_5958_p2;
wire   [0:0] xor_ln896_580_fu_5964_p2;
wire   [0:0] overflow_336_fu_5946_p2;
wire   [0:0] underflow_336_fu_5970_p2;
wire   [0:0] or_ln346_174_fu_5983_p2;
wire   [31:0] select_ln346_257_fu_5975_p3;
wire  signed [31:0] sext_ln856_165_fu_5860_p1;
wire   [19:0] zext_ln377_175_fu_6000_p1;
wire  signed [19:0] sext_ln823_166_fu_5997_p1;
wire  signed [19:0] p_Val2_852_fu_6003_p2;
wire   [0:0] p_Result_853_fu_6013_p3;
wire   [0:0] xor_ln896_514_fu_6021_p2;
wire   [0:0] xor_ln888_349_fu_6032_p2;
wire   [0:0] or_ln888_175_fu_6037_p2;
wire   [0:0] tmp_1377_fu_6048_p3;
wire   [0:0] xor_ln890_173_fu_6056_p2;
wire   [0:0] or_ln890_175_fu_6062_p2;
wire   [0:0] carry_350_fu_6027_p2;
wire   [0:0] deleted_zeros_172_fu_6043_p2;
wire   [0:0] xor_ln895_514_fu_6078_p2;
wire   [0:0] or_ln895_175_fu_6084_p2;
wire   [0:0] xor_ln895_515_fu_6090_p2;
wire   [0:0] deleted_ones_337_fu_6068_p2;
wire   [0:0] xor_ln896_515_fu_6101_p2;
wire   [0:0] and_ln891_175_fu_6073_p2;
wire   [0:0] or_ln896_175_fu_6107_p2;
wire   [0:0] xor_ln896_581_fu_6113_p2;
wire   [0:0] overflow_337_fu_6095_p2;
wire   [0:0] underflow_337_fu_6119_p2;
wire   [0:0] or_ln346_175_fu_6132_p2;
wire   [31:0] select_ln346_258_fu_6124_p3;
wire  signed [31:0] sext_ln856_166_fu_6009_p1;
wire   [30:0] zext_ln377_176_fu_6149_p1;
wire  signed [30:0] sext_ln823_167_fu_6146_p1;
wire  signed [30:0] p_Val2_855_fu_6152_p2;
wire   [0:0] p_Result_856_fu_6162_p3;
wire   [0:0] xor_ln896_516_fu_6170_p2;
wire   [0:0] xor_ln888_351_fu_6181_p2;
wire   [0:0] or_ln888_176_fu_6186_p2;
wire   [0:0] tmp_1383_fu_6197_p3;
wire   [0:0] xor_ln890_174_fu_6205_p2;
wire   [0:0] or_ln890_176_fu_6211_p2;
wire   [0:0] carry_352_fu_6176_p2;
wire   [0:0] deleted_zeros_173_fu_6192_p2;
wire   [0:0] xor_ln895_516_fu_6227_p2;
wire   [0:0] or_ln895_176_fu_6233_p2;
wire   [0:0] xor_ln895_517_fu_6239_p2;
wire   [0:0] deleted_ones_338_fu_6217_p2;
wire   [0:0] xor_ln896_517_fu_6250_p2;
wire   [0:0] and_ln891_176_fu_6222_p2;
wire   [0:0] or_ln896_176_fu_6256_p2;
wire   [0:0] xor_ln896_582_fu_6262_p2;
wire   [0:0] overflow_338_fu_6244_p2;
wire   [0:0] underflow_338_fu_6268_p2;
wire   [0:0] or_ln346_176_fu_6281_p2;
wire   [31:0] select_ln346_259_fu_6273_p3;
wire  signed [31:0] sext_ln856_167_fu_6158_p1;
wire   [30:0] zext_ln377_177_fu_6298_p1;
wire  signed [30:0] sext_ln823_168_fu_6295_p1;
wire  signed [30:0] p_Val2_858_fu_6301_p2;
wire   [0:0] p_Result_859_fu_6311_p3;
wire   [0:0] xor_ln896_518_fu_6319_p2;
wire   [0:0] xor_ln888_353_fu_6330_p2;
wire   [0:0] or_ln888_177_fu_6335_p2;
wire   [0:0] tmp_1389_fu_6346_p3;
wire   [0:0] xor_ln890_175_fu_6354_p2;
wire   [0:0] or_ln890_177_fu_6360_p2;
wire   [0:0] carry_354_fu_6325_p2;
wire   [0:0] deleted_zeros_174_fu_6341_p2;
wire   [0:0] xor_ln895_518_fu_6376_p2;
wire   [0:0] or_ln895_177_fu_6382_p2;
wire   [0:0] xor_ln895_519_fu_6388_p2;
wire   [0:0] deleted_ones_339_fu_6366_p2;
wire   [0:0] xor_ln896_519_fu_6399_p2;
wire   [0:0] and_ln891_177_fu_6371_p2;
wire   [0:0] or_ln896_177_fu_6405_p2;
wire   [0:0] xor_ln896_583_fu_6411_p2;
wire   [0:0] overflow_339_fu_6393_p2;
wire   [0:0] underflow_339_fu_6417_p2;
wire   [0:0] or_ln346_177_fu_6430_p2;
wire   [31:0] select_ln346_260_fu_6422_p3;
wire  signed [31:0] sext_ln856_168_fu_6307_p1;
wire  signed [31:0] rhs_fu_4099_p3;
wire  signed [32:0] sext_ln813_fu_6806_p1;
wire   [32:0] ret_V_fu_6810_p2;
wire   [31:0] p_Val2_887_fu_6824_p2;
wire   [0:0] p_Result_887_fu_6816_p3;
wire   [0:0] p_Result_888_fu_6830_p3;
wire   [0:0] xor_ln895_538_fu_6838_p2;
wire   [0:0] xor_ln896_538_fu_6850_p2;
wire   [0:0] xor_ln302_fu_6862_p2;
wire   [0:0] overflow_349_fu_6844_p2;
wire   [0:0] xor_ln302_323_fu_6868_p2;
wire   [0:0] underflow_349_fu_6856_p2;
wire   [0:0] or_ln302_fu_6874_p2;
wire   [31:0] select_ln302_fu_6880_p3;
wire   [31:0] select_ln350_fu_6888_p3;
wire  signed [31:0] rhs_161_fu_4224_p3;
wire  signed [32:0] sext_ln813_305_fu_6904_p1;
wire   [32:0] ret_V_161_fu_6908_p2;
wire   [31:0] p_Val2_889_fu_6922_p2;
wire   [0:0] p_Result_889_fu_6914_p3;
wire   [0:0] p_Result_890_fu_6928_p3;
wire   [0:0] xor_ln895_539_fu_6936_p2;
wire   [0:0] xor_ln896_539_fu_6948_p2;
wire   [0:0] xor_ln302_324_fu_6960_p2;
wire   [0:0] overflow_350_fu_6942_p2;
wire   [0:0] xor_ln302_325_fu_6966_p2;
wire   [0:0] underflow_350_fu_6954_p2;
wire   [0:0] or_ln302_161_fu_6972_p2;
wire   [31:0] select_ln302_324_fu_6978_p3;
wire   [31:0] select_ln350_161_fu_6986_p3;
wire  signed [31:0] rhs_162_fu_4346_p3;
wire  signed [32:0] sext_ln813_306_fu_7002_p1;
wire   [32:0] ret_V_162_fu_7006_p2;
wire   [31:0] p_Val2_891_fu_7020_p2;
wire   [0:0] p_Result_891_fu_7012_p3;
wire   [0:0] p_Result_892_fu_7026_p3;
wire   [0:0] xor_ln895_540_fu_7034_p2;
wire   [0:0] xor_ln896_540_fu_7046_p2;
wire   [0:0] xor_ln302_326_fu_7058_p2;
wire   [0:0] overflow_351_fu_7040_p2;
wire   [0:0] xor_ln302_327_fu_7064_p2;
wire   [0:0] underflow_351_fu_7052_p2;
wire   [0:0] or_ln302_162_fu_7070_p2;
wire   [31:0] select_ln302_326_fu_7076_p3;
wire   [31:0] select_ln350_162_fu_7084_p3;
wire  signed [31:0] rhs_163_fu_4470_p3;
wire  signed [32:0] sext_ln813_307_fu_7100_p1;
wire   [32:0] ret_V_163_fu_7104_p2;
wire   [31:0] p_Val2_893_fu_7118_p2;
wire   [0:0] p_Result_893_fu_7110_p3;
wire   [0:0] p_Result_894_fu_7124_p3;
wire   [0:0] xor_ln895_541_fu_7132_p2;
wire   [0:0] xor_ln896_541_fu_7144_p2;
wire   [0:0] xor_ln302_328_fu_7156_p2;
wire   [0:0] overflow_352_fu_7138_p2;
wire   [0:0] xor_ln302_329_fu_7162_p2;
wire   [0:0] underflow_352_fu_7150_p2;
wire   [0:0] or_ln302_163_fu_7168_p2;
wire   [31:0] select_ln302_328_fu_7174_p3;
wire   [31:0] select_ln350_163_fu_7182_p3;
wire  signed [31:0] rhs_164_fu_4595_p3;
wire  signed [32:0] sext_ln813_308_fu_7198_p1;
wire   [32:0] ret_V_164_fu_7202_p2;
wire   [31:0] p_Val2_895_fu_7216_p2;
wire   [0:0] p_Result_895_fu_7208_p3;
wire   [0:0] p_Result_896_fu_7222_p3;
wire   [0:0] xor_ln895_542_fu_7230_p2;
wire   [0:0] xor_ln896_542_fu_7242_p2;
wire   [0:0] xor_ln302_330_fu_7254_p2;
wire   [0:0] overflow_353_fu_7236_p2;
wire   [0:0] xor_ln302_331_fu_7260_p2;
wire   [0:0] underflow_353_fu_7248_p2;
wire   [0:0] or_ln302_164_fu_7266_p2;
wire   [31:0] select_ln302_330_fu_7272_p3;
wire   [31:0] select_ln350_164_fu_7280_p3;
wire  signed [31:0] rhs_165_fu_4720_p3;
wire  signed [32:0] sext_ln813_309_fu_7296_p1;
wire   [32:0] ret_V_165_fu_7300_p2;
wire   [31:0] p_Val2_897_fu_7314_p2;
wire   [0:0] p_Result_897_fu_7306_p3;
wire   [0:0] p_Result_898_fu_7320_p3;
wire   [0:0] xor_ln895_543_fu_7328_p2;
wire   [0:0] xor_ln896_543_fu_7340_p2;
wire   [0:0] xor_ln302_332_fu_7352_p2;
wire   [0:0] overflow_354_fu_7334_p2;
wire   [0:0] xor_ln302_333_fu_7358_p2;
wire   [0:0] underflow_354_fu_7346_p2;
wire   [0:0] or_ln302_165_fu_7364_p2;
wire   [31:0] select_ln302_332_fu_7370_p3;
wire   [31:0] select_ln350_165_fu_7378_p3;
wire  signed [31:0] rhs_166_fu_4845_p3;
wire  signed [32:0] sext_ln813_310_fu_7394_p1;
wire   [32:0] ret_V_166_fu_7398_p2;
wire   [31:0] p_Val2_899_fu_7412_p2;
wire   [0:0] p_Result_899_fu_7404_p3;
wire   [0:0] p_Result_900_fu_7418_p3;
wire   [0:0] xor_ln895_544_fu_7426_p2;
wire   [0:0] xor_ln896_544_fu_7438_p2;
wire   [0:0] xor_ln302_334_fu_7450_p2;
wire   [0:0] overflow_355_fu_7432_p2;
wire   [0:0] xor_ln302_335_fu_7456_p2;
wire   [0:0] underflow_355_fu_7444_p2;
wire   [0:0] or_ln302_166_fu_7462_p2;
wire   [31:0] select_ln302_334_fu_7468_p3;
wire   [31:0] select_ln350_166_fu_7476_p3;
wire  signed [31:0] rhs_167_fu_4970_p3;
wire  signed [32:0] sext_ln813_311_fu_7492_p1;
wire   [32:0] ret_V_167_fu_7496_p2;
wire   [31:0] p_Val2_901_fu_7510_p2;
wire   [0:0] p_Result_901_fu_7502_p3;
wire   [0:0] p_Result_902_fu_7516_p3;
wire   [0:0] xor_ln895_545_fu_7524_p2;
wire   [0:0] xor_ln896_545_fu_7536_p2;
wire   [0:0] xor_ln302_336_fu_7548_p2;
wire   [0:0] overflow_356_fu_7530_p2;
wire   [0:0] xor_ln302_337_fu_7554_p2;
wire   [0:0] underflow_356_fu_7542_p2;
wire   [0:0] or_ln302_167_fu_7560_p2;
wire   [31:0] select_ln302_336_fu_7566_p3;
wire   [31:0] select_ln350_167_fu_7574_p3;
wire  signed [31:0] rhs_168_fu_5095_p3;
wire  signed [32:0] sext_ln813_312_fu_7590_p1;
wire   [32:0] ret_V_168_fu_7594_p2;
wire   [31:0] p_Val2_903_fu_7608_p2;
wire   [0:0] p_Result_903_fu_7600_p3;
wire   [0:0] p_Result_904_fu_7614_p3;
wire   [0:0] xor_ln895_546_fu_7622_p2;
wire   [0:0] xor_ln896_546_fu_7634_p2;
wire   [0:0] xor_ln302_338_fu_7646_p2;
wire   [0:0] overflow_357_fu_7628_p2;
wire   [0:0] xor_ln302_339_fu_7652_p2;
wire   [0:0] underflow_357_fu_7640_p2;
wire   [0:0] or_ln302_168_fu_7658_p2;
wire   [31:0] select_ln302_338_fu_7664_p3;
wire   [31:0] select_ln350_168_fu_7672_p3;
wire  signed [31:0] lhs_fu_6896_p3;
wire  signed [31:0] rhs_169_fu_5244_p3;
wire  signed [32:0] sext_ln813_314_fu_7692_p1;
wire  signed [32:0] sext_ln813_313_fu_7688_p1;
wire   [32:0] ret_V_169_fu_7696_p2;
wire   [31:0] p_Val2_905_fu_7710_p2;
wire   [0:0] p_Result_905_fu_7702_p3;
wire   [0:0] p_Result_906_fu_7716_p3;
wire   [0:0] xor_ln895_547_fu_7724_p2;
wire   [0:0] xor_ln896_547_fu_7736_p2;
wire   [0:0] xor_ln302_340_fu_7748_p2;
wire   [0:0] overflow_358_fu_7730_p2;
wire   [0:0] xor_ln302_341_fu_7754_p2;
wire   [0:0] underflow_358_fu_7742_p2;
wire   [0:0] or_ln302_169_fu_7760_p2;
wire   [31:0] select_ln302_340_fu_7766_p3;
wire   [31:0] select_ln350_169_fu_7774_p3;
wire  signed [31:0] lhs_143_fu_6994_p3;
wire  signed [31:0] rhs_170_fu_5393_p3;
wire  signed [32:0] sext_ln813_316_fu_7794_p1;
wire  signed [32:0] sext_ln813_315_fu_7790_p1;
wire   [32:0] ret_V_170_fu_7798_p2;
wire   [31:0] p_Val2_907_fu_7812_p2;
wire   [0:0] p_Result_907_fu_7804_p3;
wire   [0:0] p_Result_908_fu_7818_p3;
wire   [0:0] xor_ln895_548_fu_7826_p2;
wire   [0:0] xor_ln896_548_fu_7838_p2;
wire   [0:0] xor_ln302_342_fu_7850_p2;
wire   [0:0] overflow_359_fu_7832_p2;
wire   [0:0] xor_ln302_343_fu_7856_p2;
wire   [0:0] underflow_359_fu_7844_p2;
wire   [0:0] or_ln302_170_fu_7862_p2;
wire   [31:0] select_ln302_342_fu_7868_p3;
wire   [31:0] select_ln350_170_fu_7876_p3;
wire  signed [31:0] lhs_144_fu_7092_p3;
wire  signed [31:0] rhs_171_fu_5542_p3;
wire  signed [32:0] sext_ln813_318_fu_7896_p1;
wire  signed [32:0] sext_ln813_317_fu_7892_p1;
wire   [32:0] ret_V_171_fu_7900_p2;
wire   [31:0] p_Val2_909_fu_7914_p2;
wire   [0:0] p_Result_909_fu_7906_p3;
wire   [0:0] p_Result_910_fu_7920_p3;
wire   [0:0] xor_ln895_549_fu_7928_p2;
wire   [0:0] xor_ln896_549_fu_7940_p2;
wire   [0:0] xor_ln302_344_fu_7952_p2;
wire   [0:0] overflow_360_fu_7934_p2;
wire   [0:0] xor_ln302_345_fu_7958_p2;
wire   [0:0] underflow_360_fu_7946_p2;
wire   [0:0] or_ln302_171_fu_7964_p2;
wire   [31:0] select_ln302_344_fu_7970_p3;
wire   [31:0] select_ln350_171_fu_7978_p3;
wire  signed [31:0] lhs_145_fu_7190_p3;
wire  signed [31:0] rhs_172_fu_5691_p3;
wire  signed [32:0] sext_ln813_320_fu_7998_p1;
wire  signed [32:0] sext_ln813_319_fu_7994_p1;
wire   [32:0] ret_V_172_fu_8002_p2;
wire   [31:0] p_Val2_911_fu_8016_p2;
wire   [0:0] p_Result_911_fu_8008_p3;
wire   [0:0] p_Result_912_fu_8022_p3;
wire   [0:0] xor_ln895_550_fu_8030_p2;
wire   [0:0] xor_ln896_550_fu_8042_p2;
wire   [0:0] xor_ln302_346_fu_8054_p2;
wire   [0:0] overflow_361_fu_8036_p2;
wire   [0:0] xor_ln302_347_fu_8060_p2;
wire   [0:0] underflow_361_fu_8048_p2;
wire   [0:0] or_ln302_172_fu_8066_p2;
wire   [31:0] select_ln302_346_fu_8072_p3;
wire   [31:0] select_ln350_172_fu_8080_p3;
wire  signed [31:0] lhs_146_fu_7288_p3;
wire  signed [31:0] rhs_173_fu_5840_p3;
wire  signed [32:0] sext_ln813_322_fu_8100_p1;
wire  signed [32:0] sext_ln813_321_fu_8096_p1;
wire   [32:0] ret_V_173_fu_8104_p2;
wire   [31:0] p_Val2_913_fu_8118_p2;
wire   [0:0] p_Result_913_fu_8110_p3;
wire   [0:0] p_Result_914_fu_8124_p3;
wire   [0:0] xor_ln895_551_fu_8132_p2;
wire   [0:0] xor_ln896_551_fu_8144_p2;
wire   [0:0] xor_ln302_348_fu_8156_p2;
wire   [0:0] overflow_362_fu_8138_p2;
wire   [0:0] xor_ln302_349_fu_8162_p2;
wire   [0:0] underflow_362_fu_8150_p2;
wire   [0:0] or_ln302_173_fu_8168_p2;
wire   [31:0] select_ln302_348_fu_8174_p3;
wire   [31:0] select_ln350_173_fu_8182_p3;
wire  signed [31:0] lhs_147_fu_7386_p3;
wire  signed [31:0] rhs_174_fu_5989_p3;
wire  signed [32:0] sext_ln813_324_fu_8202_p1;
wire  signed [32:0] sext_ln813_323_fu_8198_p1;
wire   [32:0] ret_V_174_fu_8206_p2;
wire   [31:0] p_Val2_915_fu_8220_p2;
wire   [0:0] p_Result_915_fu_8212_p3;
wire   [0:0] p_Result_916_fu_8226_p3;
wire   [0:0] xor_ln895_552_fu_8234_p2;
wire   [0:0] xor_ln896_552_fu_8246_p2;
wire   [0:0] xor_ln302_350_fu_8258_p2;
wire   [0:0] overflow_363_fu_8240_p2;
wire   [0:0] xor_ln302_351_fu_8264_p2;
wire   [0:0] underflow_363_fu_8252_p2;
wire   [0:0] or_ln302_174_fu_8270_p2;
wire   [31:0] select_ln302_350_fu_8276_p3;
wire   [31:0] select_ln350_174_fu_8284_p3;
wire  signed [31:0] lhs_148_fu_7484_p3;
wire  signed [31:0] rhs_175_fu_6138_p3;
wire  signed [32:0] sext_ln813_326_fu_8304_p1;
wire  signed [32:0] sext_ln813_325_fu_8300_p1;
wire   [32:0] ret_V_175_fu_8308_p2;
wire   [31:0] p_Val2_917_fu_8322_p2;
wire   [0:0] p_Result_917_fu_8314_p3;
wire   [0:0] p_Result_918_fu_8328_p3;
wire   [0:0] xor_ln895_553_fu_8336_p2;
wire   [0:0] xor_ln896_553_fu_8348_p2;
wire   [0:0] xor_ln302_352_fu_8360_p2;
wire   [0:0] overflow_364_fu_8342_p2;
wire   [0:0] xor_ln302_353_fu_8366_p2;
wire   [0:0] underflow_364_fu_8354_p2;
wire   [0:0] or_ln302_175_fu_8372_p2;
wire   [31:0] select_ln302_352_fu_8378_p3;
wire   [31:0] select_ln350_175_fu_8386_p3;
wire  signed [31:0] lhs_149_fu_7582_p3;
wire  signed [31:0] rhs_176_fu_6287_p3;
wire  signed [32:0] sext_ln813_328_fu_8406_p1;
wire  signed [32:0] sext_ln813_327_fu_8402_p1;
wire   [32:0] ret_V_176_fu_8410_p2;
wire   [31:0] p_Val2_919_fu_8424_p2;
wire   [0:0] p_Result_919_fu_8416_p3;
wire   [0:0] p_Result_920_fu_8430_p3;
wire   [0:0] xor_ln895_554_fu_8438_p2;
wire   [0:0] xor_ln896_554_fu_8450_p2;
wire   [0:0] xor_ln302_354_fu_8462_p2;
wire   [0:0] overflow_365_fu_8444_p2;
wire   [0:0] xor_ln302_355_fu_8468_p2;
wire   [0:0] underflow_365_fu_8456_p2;
wire   [0:0] or_ln302_176_fu_8474_p2;
wire   [31:0] select_ln302_354_fu_8480_p3;
wire   [31:0] select_ln350_176_fu_8488_p3;
wire  signed [31:0] lhs_150_fu_7680_p3;
wire  signed [31:0] rhs_177_fu_6436_p3;
wire  signed [32:0] sext_ln813_330_fu_8508_p1;
wire  signed [32:0] sext_ln813_329_fu_8504_p1;
wire   [32:0] ret_V_177_fu_8512_p2;
wire   [31:0] p_Val2_921_fu_8526_p2;
wire   [0:0] p_Result_921_fu_8518_p3;
wire   [0:0] p_Result_922_fu_8532_p3;
wire   [0:0] xor_ln895_555_fu_8540_p2;
wire   [0:0] xor_ln896_555_fu_8552_p2;
wire   [0:0] xor_ln302_356_fu_8564_p2;
wire   [0:0] overflow_366_fu_8546_p2;
wire   [0:0] xor_ln302_357_fu_8570_p2;
wire   [0:0] underflow_366_fu_8558_p2;
wire   [0:0] or_ln302_177_fu_8576_p2;
wire   [31:0] select_ln302_356_fu_8582_p3;
wire   [31:0] select_ln350_177_fu_8590_p3;
wire   [19:0] zext_ln377_178_fu_8609_p1;
wire  signed [19:0] sext_ln823_169_fu_8606_p1;
wire  signed [19:0] p_Val2_861_fu_8612_p2;
wire   [0:0] p_Result_862_fu_8622_p3;
wire   [0:0] xor_ln896_520_fu_8630_p2;
wire   [0:0] xor_ln888_355_fu_8641_p2;
wire   [0:0] or_ln888_178_fu_8646_p2;
wire   [0:0] tmp_1395_fu_8657_p3;
wire   [0:0] xor_ln890_176_fu_8665_p2;
wire   [0:0] or_ln890_178_fu_8671_p2;
wire   [0:0] carry_356_fu_8636_p2;
wire   [0:0] deleted_zeros_175_fu_8652_p2;
wire   [0:0] xor_ln895_520_fu_8687_p2;
wire   [0:0] or_ln895_178_fu_8693_p2;
wire   [0:0] xor_ln895_521_fu_8699_p2;
wire   [0:0] deleted_ones_340_fu_8677_p2;
wire   [0:0] xor_ln896_521_fu_8710_p2;
wire   [0:0] and_ln891_178_fu_8682_p2;
wire   [0:0] or_ln896_178_fu_8716_p2;
wire   [0:0] xor_ln896_584_fu_8722_p2;
wire   [0:0] overflow_340_fu_8704_p2;
wire   [0:0] underflow_340_fu_8728_p2;
wire   [0:0] or_ln346_178_fu_8741_p2;
wire   [31:0] select_ln346_261_fu_8733_p3;
wire  signed [31:0] sext_ln856_169_fu_8618_p1;
wire   [18:0] zext_ln377_179_fu_8758_p1;
wire  signed [18:0] sext_ln823_170_fu_8755_p1;
wire  signed [18:0] p_Val2_864_fu_8761_p2;
wire   [0:0] p_Result_865_fu_8771_p3;
wire   [0:0] xor_ln896_522_fu_8779_p2;
wire   [0:0] xor_ln888_357_fu_8790_p2;
wire   [0:0] or_ln888_179_fu_8795_p2;
wire   [0:0] tmp_1401_fu_8806_p3;
wire   [0:0] xor_ln890_177_fu_8814_p2;
wire   [0:0] or_ln890_179_fu_8820_p2;
wire   [0:0] carry_358_fu_8785_p2;
wire   [0:0] deleted_zeros_176_fu_8801_p2;
wire   [0:0] xor_ln895_522_fu_8836_p2;
wire   [0:0] or_ln895_179_fu_8842_p2;
wire   [0:0] xor_ln895_523_fu_8848_p2;
wire   [0:0] deleted_ones_341_fu_8826_p2;
wire   [0:0] xor_ln896_523_fu_8859_p2;
wire   [0:0] and_ln891_179_fu_8831_p2;
wire   [0:0] or_ln896_179_fu_8865_p2;
wire   [0:0] xor_ln896_585_fu_8871_p2;
wire   [0:0] overflow_341_fu_8853_p2;
wire   [0:0] underflow_341_fu_8877_p2;
wire   [0:0] or_ln346_179_fu_8890_p2;
wire   [31:0] select_ln346_262_fu_8882_p3;
wire  signed [31:0] sext_ln856_170_fu_8767_p1;
wire   [20:0] zext_ln377_180_fu_8907_p1;
wire  signed [20:0] sext_ln823_171_fu_8904_p1;
wire  signed [20:0] p_Val2_867_fu_8910_p2;
wire   [0:0] p_Result_868_fu_8920_p3;
wire   [0:0] xor_ln896_524_fu_8928_p2;
wire   [0:0] xor_ln888_359_fu_8939_p2;
wire   [0:0] or_ln888_180_fu_8944_p2;
wire   [0:0] tmp_1407_fu_8955_p3;
wire   [0:0] xor_ln890_178_fu_8963_p2;
wire   [0:0] or_ln890_180_fu_8969_p2;
wire   [0:0] carry_360_fu_8934_p2;
wire   [0:0] deleted_zeros_177_fu_8950_p2;
wire   [0:0] xor_ln895_524_fu_8985_p2;
wire   [0:0] or_ln895_180_fu_8991_p2;
wire   [0:0] xor_ln895_525_fu_8997_p2;
wire   [0:0] deleted_ones_342_fu_8975_p2;
wire   [0:0] xor_ln896_525_fu_9008_p2;
wire   [0:0] and_ln891_180_fu_8980_p2;
wire   [0:0] or_ln896_180_fu_9014_p2;
wire   [0:0] xor_ln896_586_fu_9020_p2;
wire   [0:0] overflow_342_fu_9002_p2;
wire   [0:0] underflow_342_fu_9026_p2;
wire   [0:0] or_ln346_180_fu_9039_p2;
wire   [31:0] select_ln346_263_fu_9031_p3;
wire  signed [31:0] sext_ln856_171_fu_8916_p1;
wire   [21:0] zext_ln377_181_fu_9056_p1;
wire  signed [21:0] sext_ln823_172_fu_9053_p1;
wire  signed [21:0] p_Val2_870_fu_9059_p2;
wire   [0:0] p_Result_871_fu_9069_p3;
wire   [0:0] xor_ln896_526_fu_9077_p2;
wire   [0:0] xor_ln888_361_fu_9088_p2;
wire   [0:0] or_ln888_181_fu_9093_p2;
wire   [0:0] tmp_1413_fu_9104_p3;
wire   [0:0] xor_ln890_179_fu_9112_p2;
wire   [0:0] or_ln890_181_fu_9118_p2;
wire   [0:0] carry_362_fu_9083_p2;
wire   [0:0] deleted_zeros_178_fu_9099_p2;
wire   [0:0] xor_ln895_526_fu_9134_p2;
wire   [0:0] or_ln895_181_fu_9140_p2;
wire   [0:0] xor_ln895_527_fu_9146_p2;
wire   [0:0] deleted_ones_343_fu_9124_p2;
wire   [0:0] xor_ln896_527_fu_9157_p2;
wire   [0:0] and_ln891_181_fu_9129_p2;
wire   [0:0] or_ln896_181_fu_9163_p2;
wire   [0:0] xor_ln896_587_fu_9169_p2;
wire   [0:0] overflow_343_fu_9151_p2;
wire   [0:0] underflow_343_fu_9175_p2;
wire   [0:0] or_ln346_181_fu_9188_p2;
wire   [31:0] select_ln346_264_fu_9180_p3;
wire  signed [31:0] sext_ln856_172_fu_9065_p1;
wire   [30:0] zext_ln377_182_fu_9205_p1;
wire  signed [30:0] sext_ln823_173_fu_9202_p1;
wire  signed [30:0] p_Val2_873_fu_9208_p2;
wire   [0:0] p_Result_874_fu_9218_p3;
wire   [0:0] xor_ln896_528_fu_9226_p2;
wire   [0:0] xor_ln888_363_fu_9237_p2;
wire   [0:0] or_ln888_182_fu_9242_p2;
wire   [0:0] tmp_1419_fu_9253_p3;
wire   [0:0] xor_ln890_180_fu_9261_p2;
wire   [0:0] or_ln890_182_fu_9267_p2;
wire   [0:0] carry_364_fu_9232_p2;
wire   [0:0] deleted_zeros_179_fu_9248_p2;
wire   [0:0] xor_ln895_528_fu_9283_p2;
wire   [0:0] or_ln895_182_fu_9289_p2;
wire   [0:0] xor_ln895_529_fu_9295_p2;
wire   [0:0] deleted_ones_344_fu_9273_p2;
wire   [0:0] xor_ln896_529_fu_9306_p2;
wire   [0:0] and_ln891_182_fu_9278_p2;
wire   [0:0] or_ln896_182_fu_9312_p2;
wire   [0:0] xor_ln896_588_fu_9318_p2;
wire   [0:0] overflow_344_fu_9300_p2;
wire   [0:0] underflow_344_fu_9324_p2;
wire   [0:0] or_ln346_182_fu_9337_p2;
wire   [31:0] select_ln346_265_fu_9329_p3;
wire  signed [31:0] sext_ln856_173_fu_9214_p1;
wire   [31:0] select_ln346_266_fu_9354_p3;
wire  signed [31:0] sext_ln856_174_fu_9351_p1;
wire   [17:0] zext_ln377_184_fu_9371_p1;
wire  signed [17:0] sext_ln823_175_fu_9368_p1;
wire  signed [17:0] p_Val2_879_fu_9374_p2;
wire   [0:0] p_Result_880_fu_9384_p3;
wire   [0:0] xor_ln896_532_fu_9392_p2;
wire   [0:0] xor_ln888_367_fu_9403_p2;
wire   [0:0] or_ln888_184_fu_9408_p2;
wire   [0:0] tmp_1431_fu_9419_p3;
wire   [0:0] xor_ln890_182_fu_9427_p2;
wire   [0:0] or_ln890_184_fu_9433_p2;
wire   [0:0] carry_368_fu_9398_p2;
wire   [0:0] deleted_zeros_181_fu_9414_p2;
wire   [0:0] xor_ln895_532_fu_9449_p2;
wire   [0:0] or_ln895_184_fu_9455_p2;
wire   [0:0] xor_ln895_533_fu_9461_p2;
wire   [0:0] deleted_ones_346_fu_9439_p2;
wire   [0:0] xor_ln896_533_fu_9472_p2;
wire   [0:0] and_ln891_184_fu_9444_p2;
wire   [0:0] or_ln896_184_fu_9478_p2;
wire   [0:0] xor_ln896_590_fu_9484_p2;
wire   [0:0] overflow_346_fu_9466_p2;
wire   [0:0] underflow_346_fu_9490_p2;
wire   [0:0] or_ln346_184_fu_9503_p2;
wire   [31:0] select_ln346_267_fu_9495_p3;
wire  signed [31:0] sext_ln856_175_fu_9380_p1;
wire   [30:0] zext_ln377_185_fu_9520_p1;
wire  signed [30:0] sext_ln823_176_fu_9517_p1;
wire  signed [30:0] p_Val2_882_fu_9523_p2;
wire   [0:0] p_Result_883_fu_9533_p3;
wire   [0:0] xor_ln896_534_fu_9541_p2;
wire   [0:0] xor_ln888_369_fu_9552_p2;
wire   [0:0] or_ln888_185_fu_9557_p2;
wire   [0:0] tmp_1437_fu_9568_p3;
wire   [0:0] xor_ln890_183_fu_9576_p2;
wire   [0:0] or_ln890_185_fu_9582_p2;
wire   [0:0] carry_370_fu_9547_p2;
wire   [0:0] deleted_zeros_182_fu_9563_p2;
wire   [0:0] xor_ln895_534_fu_9598_p2;
wire   [0:0] or_ln895_185_fu_9604_p2;
wire   [0:0] xor_ln895_535_fu_9610_p2;
wire   [0:0] deleted_ones_347_fu_9588_p2;
wire   [0:0] xor_ln896_535_fu_9621_p2;
wire   [0:0] and_ln891_185_fu_9593_p2;
wire   [0:0] or_ln896_185_fu_9627_p2;
wire   [0:0] xor_ln896_591_fu_9633_p2;
wire   [0:0] overflow_347_fu_9615_p2;
wire   [0:0] underflow_347_fu_9639_p2;
wire   [0:0] or_ln346_185_fu_9652_p2;
wire   [31:0] select_ln346_268_fu_9644_p3;
wire  signed [31:0] sext_ln856_176_fu_9529_p1;
wire   [30:0] zext_ln377_186_fu_9669_p1;
wire  signed [30:0] sext_ln823_177_fu_9666_p1;
wire  signed [30:0] p_Val2_885_fu_9672_p2;
wire   [0:0] p_Result_886_fu_9682_p3;
wire   [0:0] xor_ln896_536_fu_9690_p2;
wire   [0:0] xor_ln888_371_fu_9701_p2;
wire   [0:0] or_ln888_186_fu_9706_p2;
wire   [0:0] tmp_1443_fu_9717_p3;
wire   [0:0] xor_ln890_184_fu_9725_p2;
wire   [0:0] or_ln890_186_fu_9731_p2;
wire   [0:0] carry_372_fu_9696_p2;
wire   [0:0] deleted_zeros_183_fu_9712_p2;
wire   [0:0] xor_ln895_536_fu_9747_p2;
wire   [0:0] or_ln895_186_fu_9753_p2;
wire   [0:0] xor_ln895_537_fu_9759_p2;
wire   [0:0] deleted_ones_348_fu_9737_p2;
wire   [0:0] xor_ln896_537_fu_9770_p2;
wire   [0:0] and_ln891_186_fu_9742_p2;
wire   [0:0] or_ln896_186_fu_9776_p2;
wire   [0:0] xor_ln896_592_fu_9782_p2;
wire   [0:0] overflow_348_fu_9764_p2;
wire   [0:0] underflow_348_fu_9788_p2;
wire   [0:0] or_ln346_186_fu_9801_p2;
wire   [31:0] select_ln346_269_fu_9793_p3;
wire  signed [31:0] sext_ln856_177_fu_9678_p1;
wire  signed [31:0] rhs_178_fu_8747_p3;
wire  signed [32:0] sext_ln813_332_fu_9818_p1;
wire  signed [32:0] sext_ln813_331_fu_9815_p1;
wire   [32:0] ret_V_178_fu_9822_p2;
wire   [31:0] p_Val2_923_fu_9836_p2;
wire   [0:0] p_Result_923_fu_9828_p3;
wire   [0:0] p_Result_924_fu_9841_p3;
wire   [0:0] xor_ln895_556_fu_9849_p2;
wire   [0:0] xor_ln896_556_fu_9861_p2;
wire   [0:0] xor_ln302_358_fu_9873_p2;
wire   [0:0] overflow_367_fu_9855_p2;
wire   [0:0] xor_ln302_359_fu_9879_p2;
wire   [0:0] underflow_367_fu_9867_p2;
wire   [0:0] or_ln302_178_fu_9885_p2;
wire   [31:0] select_ln302_358_fu_9891_p3;
wire   [31:0] select_ln350_178_fu_9899_p3;
wire  signed [31:0] rhs_179_fu_8896_p3;
wire  signed [32:0] sext_ln813_334_fu_9918_p1;
wire  signed [32:0] sext_ln813_333_fu_9915_p1;
wire   [32:0] ret_V_179_fu_9922_p2;
wire   [31:0] p_Val2_925_fu_9936_p2;
wire   [0:0] p_Result_925_fu_9928_p3;
wire   [0:0] p_Result_926_fu_9941_p3;
wire   [0:0] xor_ln895_557_fu_9949_p2;
wire   [0:0] xor_ln896_557_fu_9961_p2;
wire   [0:0] xor_ln302_360_fu_9973_p2;
wire   [0:0] overflow_368_fu_9955_p2;
wire   [0:0] xor_ln302_361_fu_9979_p2;
wire   [0:0] underflow_368_fu_9967_p2;
wire   [0:0] or_ln302_179_fu_9985_p2;
wire   [31:0] select_ln302_360_fu_9991_p3;
wire   [31:0] select_ln350_179_fu_9999_p3;
wire  signed [31:0] rhs_180_fu_9045_p3;
wire  signed [32:0] sext_ln813_336_fu_10018_p1;
wire  signed [32:0] sext_ln813_335_fu_10015_p1;
wire   [32:0] ret_V_180_fu_10022_p2;
wire   [31:0] p_Val2_927_fu_10036_p2;
wire   [0:0] p_Result_927_fu_10028_p3;
wire   [0:0] p_Result_928_fu_10041_p3;
wire   [0:0] xor_ln895_558_fu_10049_p2;
wire   [0:0] xor_ln896_558_fu_10061_p2;
wire   [0:0] xor_ln302_362_fu_10073_p2;
wire   [0:0] overflow_369_fu_10055_p2;
wire   [0:0] xor_ln302_363_fu_10079_p2;
wire   [0:0] underflow_369_fu_10067_p2;
wire   [0:0] or_ln302_180_fu_10085_p2;
wire   [31:0] select_ln302_362_fu_10091_p3;
wire   [31:0] select_ln350_180_fu_10099_p3;
wire  signed [31:0] rhs_181_fu_9194_p3;
wire  signed [32:0] sext_ln813_338_fu_10118_p1;
wire  signed [32:0] sext_ln813_337_fu_10115_p1;
wire   [32:0] ret_V_181_fu_10122_p2;
wire   [31:0] p_Val2_929_fu_10136_p2;
wire   [0:0] p_Result_929_fu_10128_p3;
wire   [0:0] p_Result_930_fu_10141_p3;
wire   [0:0] xor_ln895_559_fu_10149_p2;
wire   [0:0] xor_ln896_559_fu_10161_p2;
wire   [0:0] xor_ln302_364_fu_10173_p2;
wire   [0:0] overflow_370_fu_10155_p2;
wire   [0:0] xor_ln302_365_fu_10179_p2;
wire   [0:0] underflow_370_fu_10167_p2;
wire   [0:0] or_ln302_181_fu_10185_p2;
wire   [31:0] select_ln302_364_fu_10191_p3;
wire   [31:0] select_ln350_181_fu_10199_p3;
wire  signed [31:0] rhs_182_fu_9343_p3;
wire  signed [32:0] sext_ln813_340_fu_10218_p1;
wire  signed [32:0] sext_ln813_339_fu_10215_p1;
wire   [32:0] ret_V_182_fu_10222_p2;
wire   [31:0] p_Val2_931_fu_10236_p2;
wire   [0:0] p_Result_931_fu_10228_p3;
wire   [0:0] p_Result_932_fu_10241_p3;
wire   [0:0] xor_ln895_560_fu_10249_p2;
wire   [0:0] xor_ln896_560_fu_10261_p2;
wire   [0:0] xor_ln302_366_fu_10273_p2;
wire   [0:0] overflow_371_fu_10255_p2;
wire   [0:0] xor_ln302_367_fu_10279_p2;
wire   [0:0] underflow_371_fu_10267_p2;
wire   [0:0] or_ln302_182_fu_10285_p2;
wire   [31:0] select_ln302_366_fu_10291_p3;
wire   [31:0] select_ln350_182_fu_10299_p3;
wire  signed [31:0] rhs_183_fu_9361_p3;
wire  signed [32:0] sext_ln813_342_fu_10318_p1;
wire  signed [32:0] sext_ln813_341_fu_10315_p1;
wire   [32:0] ret_V_183_fu_10322_p2;
wire   [31:0] p_Val2_933_fu_10336_p2;
wire   [0:0] p_Result_933_fu_10328_p3;
wire   [0:0] p_Result_934_fu_10341_p3;
wire   [0:0] xor_ln895_561_fu_10349_p2;
wire   [0:0] xor_ln896_561_fu_10361_p2;
wire   [0:0] xor_ln302_368_fu_10373_p2;
wire   [0:0] overflow_372_fu_10355_p2;
wire   [0:0] xor_ln302_369_fu_10379_p2;
wire   [0:0] underflow_372_fu_10367_p2;
wire   [0:0] or_ln302_183_fu_10385_p2;
wire   [31:0] select_ln302_368_fu_10391_p3;
wire   [31:0] select_ln350_183_fu_10399_p3;
wire  signed [31:0] rhs_184_fu_9509_p3;
wire  signed [32:0] sext_ln813_344_fu_10418_p1;
wire  signed [32:0] sext_ln813_343_fu_10415_p1;
wire   [32:0] ret_V_184_fu_10422_p2;
wire   [31:0] p_Val2_935_fu_10436_p2;
wire   [0:0] p_Result_935_fu_10428_p3;
wire   [0:0] p_Result_936_fu_10441_p3;
wire   [0:0] xor_ln895_562_fu_10449_p2;
wire   [0:0] xor_ln896_562_fu_10461_p2;
wire   [0:0] xor_ln302_370_fu_10473_p2;
wire   [0:0] overflow_373_fu_10455_p2;
wire   [0:0] xor_ln302_371_fu_10479_p2;
wire   [0:0] underflow_373_fu_10467_p2;
wire   [0:0] or_ln302_184_fu_10485_p2;
wire   [31:0] select_ln302_370_fu_10491_p3;
wire   [31:0] select_ln350_184_fu_10499_p3;
wire  signed [31:0] rhs_185_fu_9658_p3;
wire  signed [32:0] sext_ln813_346_fu_10518_p1;
wire  signed [32:0] sext_ln813_345_fu_10515_p1;
wire   [32:0] ret_V_185_fu_10522_p2;
wire   [31:0] p_Val2_937_fu_10536_p2;
wire   [0:0] p_Result_937_fu_10528_p3;
wire   [0:0] p_Result_938_fu_10541_p3;
wire   [0:0] xor_ln895_563_fu_10549_p2;
wire   [0:0] xor_ln896_563_fu_10561_p2;
wire   [0:0] xor_ln302_372_fu_10573_p2;
wire   [0:0] overflow_374_fu_10555_p2;
wire   [0:0] xor_ln302_373_fu_10579_p2;
wire   [0:0] underflow_374_fu_10567_p2;
wire   [0:0] or_ln302_185_fu_10585_p2;
wire   [31:0] select_ln302_372_fu_10591_p3;
wire   [31:0] select_ln350_185_fu_10599_p3;
wire  signed [31:0] rhs_186_fu_9807_p3;
wire  signed [32:0] sext_ln813_348_fu_10618_p1;
wire  signed [32:0] sext_ln813_347_fu_10615_p1;
wire   [32:0] ret_V_186_fu_10622_p2;
wire   [31:0] p_Val2_939_fu_10636_p2;
wire   [0:0] p_Result_939_fu_10628_p3;
wire   [0:0] p_Result_940_fu_10641_p3;
wire   [0:0] xor_ln895_564_fu_10649_p2;
wire   [0:0] xor_ln896_564_fu_10661_p2;
wire   [0:0] xor_ln302_374_fu_10673_p2;
wire   [0:0] overflow_375_fu_10655_p2;
wire   [0:0] xor_ln302_375_fu_10679_p2;
wire   [0:0] underflow_375_fu_10667_p2;
wire   [0:0] or_ln302_186_fu_10685_p2;
wire   [31:0] select_ln302_374_fu_10691_p3;
wire   [31:0] select_ln350_186_fu_10699_p3;
wire   [31:0] select_ln302_359_fu_9907_p3;
wire   [31:0] select_ln302_361_fu_10007_p3;
wire   [31:0] select_ln302_363_fu_10107_p3;
wire   [31:0] select_ln302_365_fu_10207_p3;
wire   [31:0] select_ln302_367_fu_10307_p3;
wire   [31:0] select_ln302_369_fu_10407_p3;
wire   [31:0] select_ln302_371_fu_10507_p3;
wire   [31:0] select_ln302_373_fu_10607_p3;
wire   [31:0] select_ln302_375_fu_10707_p3;
reg    ap_ce_reg;
reg   [95:0] p_read_int_reg;
reg   [31:0] ap_return_0_int_reg;
reg   [31:0] ap_return_1_int_reg;
reg   [31:0] ap_return_2_int_reg;
reg   [31:0] ap_return_3_int_reg;
reg   [31:0] ap_return_4_int_reg;
reg   [31:0] ap_return_5_int_reg;
reg   [31:0] ap_return_6_int_reg;
reg   [31:0] ap_return_7_int_reg;
reg   [31:0] ap_return_8_int_reg;

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U1(
    .din0(r_V_183_fu_240_p0),
    .din1(r_V_183_fu_240_p1),
    .dout(r_V_183_fu_240_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U2(
    .din0(a_V_1_fu_3313_p4),
    .din1(r_V_189_fu_242_p1),
    .dout(r_V_189_fu_242_p2)
);

motorB_mul_32s_23s_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23s_54_1_0_U3(
    .din0(r_V_194_fu_243_p0),
    .din1(r_V_194_fu_243_p1),
    .dout(r_V_194_fu_243_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U4(
    .din0(r_V_193_fu_244_p0),
    .din1(r_V_193_fu_244_p1),
    .dout(r_V_193_fu_244_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U5(
    .din0(a_V_2_reg_11309),
    .din1(r_V_197_fu_245_p1),
    .dout(r_V_197_fu_245_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U6(
    .din0(r_V_186_fu_246_p0),
    .din1(r_V_186_fu_246_p1),
    .dout(r_V_186_fu_246_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U7(
    .din0(a_V_2_reg_11309),
    .din1(r_V_fu_247_p1),
    .dout(r_V_fu_247_p2)
);

motorB_mul_32s_23s_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23s_54_1_0_U8(
    .din0(r_V_195_fu_248_p0),
    .din1(r_V_195_fu_248_p1),
    .dout(r_V_195_fu_248_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U9(
    .din0(r_V_184_fu_249_p0),
    .din1(r_V_184_fu_249_p1),
    .dout(r_V_184_fu_249_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U10(
    .din0(r_V_192_fu_250_p0),
    .din1(r_V_192_fu_250_p1),
    .dout(r_V_192_fu_250_p2)
);

motorB_mul_32s_26ns_57_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 26 ),
    .dout_WIDTH( 57 ))
mul_32s_26ns_57_1_0_U11(
    .din0(a_V_fu_2708_p1),
    .din1(r_V_180_fu_251_p1),
    .dout(r_V_180_fu_251_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U12(
    .din0(r_V_202_fu_252_p0),
    .din1(r_V_202_fu_252_p1),
    .dout(r_V_202_fu_252_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U13(
    .din0(r_V_203_fu_253_p0),
    .din1(r_V_203_fu_253_p1),
    .dout(r_V_203_fu_253_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U14(
    .din0(r_V_178_fu_254_p0),
    .din1(r_V_178_fu_254_p1),
    .dout(r_V_178_fu_254_p2)
);

motorB_mul_32s_23s_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23s_54_1_0_U15(
    .din0(r_V_199_fu_255_p0),
    .din1(r_V_199_fu_255_p1),
    .dout(r_V_199_fu_255_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U16(
    .din0(r_V_181_fu_256_p0),
    .din1(r_V_181_fu_256_p1),
    .dout(r_V_181_fu_256_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U17(
    .din0(a_V_2_reg_11309),
    .din1(r_V_201_fu_257_p1),
    .dout(r_V_201_fu_257_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U18(
    .din0(a_V_2_reg_11309),
    .din1(r_V_196_fu_258_p1),
    .dout(r_V_196_fu_258_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U19(
    .din0(r_V_185_fu_259_p0),
    .din1(r_V_185_fu_259_p1),
    .dout(r_V_185_fu_259_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U20(
    .din0(r_V_190_fu_260_p0),
    .din1(r_V_190_fu_260_p1),
    .dout(r_V_190_fu_260_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U21(
    .din0(r_V_188_fu_261_p0),
    .din1(r_V_188_fu_261_p1),
    .dout(r_V_188_fu_261_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U22(
    .din0(r_V_179_fu_262_p0),
    .din1(r_V_179_fu_262_p1),
    .dout(r_V_179_fu_262_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U23(
    .din0(r_V_191_fu_263_p0),
    .din1(r_V_191_fu_263_p1),
    .dout(r_V_191_fu_263_p2)
);

motorB_mul_32s_15ns_47_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 47 ))
mul_32s_15ns_47_1_0_U24(
    .din0(a_V_fu_2708_p1),
    .din1(r_V_182_fu_264_p1),
    .dout(r_V_182_fu_264_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U25(
    .din0(a_V_2_reg_11309),
    .din1(r_V_198_fu_265_p1),
    .dout(r_V_198_fu_265_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U26(
    .din0(a_V_1_fu_3313_p4),
    .din1(r_V_187_fu_266_p1),
    .dout(r_V_187_fu_266_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        Range2_all_ones_159_reg_10824 <= r_V_179_fu_262_p2[32'd43];
        Range2_all_ones_160_reg_10855 <= r_V_180_fu_251_p2[32'd56];
        Range2_all_ones_161_reg_10886 <= r_V_181_fu_256_p2[32'd43];
        Range2_all_ones_162_reg_10917 <= r_V_182_fu_264_p2[32'd46];
        Range2_all_ones_163_reg_10948 <= r_V_183_fu_240_p2[32'd42];
        Range2_all_ones_164_reg_10979 <= r_V_184_fu_249_p2[32'd42];
        Range2_all_ones_165_reg_11010 <= r_V_185_fu_259_p2[32'd53];
        Range2_all_ones_166_reg_11041 <= r_V_186_fu_246_p2[32'd53];
        Range2_all_ones_167_reg_11070 <= r_V_187_fu_266_p2[32'd40];
        Range2_all_ones_168_reg_11099 <= r_V_188_fu_261_p2[32'd42];
        Range2_all_ones_169_reg_11128 <= r_V_189_fu_242_p2[32'd44];
        Range2_all_ones_170_reg_11157 <= r_V_190_fu_260_p2[32'd42];
        Range2_all_ones_171_reg_11186 <= r_V_191_fu_263_p2[32'd53];
        Range2_all_ones_172_reg_11215 <= r_V_192_fu_250_p2[32'd42];
        Range2_all_ones_173_reg_11244 <= r_V_193_fu_244_p2[32'd42];
        Range2_all_ones_174_reg_11273 <= r_V_194_fu_243_p2[32'd53];
        Range2_all_ones_175_reg_11302 <= r_V_195_fu_248_p2[32'd53];
        Range2_all_ones_176_reg_11356 <= r_V_fu_247_p2[32'd42];
        Range2_all_ones_177_reg_11385 <= r_V_196_fu_258_p2[32'd41];
        Range2_all_ones_178_reg_11414 <= r_V_197_fu_245_p2[32'd43];
        Range2_all_ones_179_reg_11443 <= r_V_198_fu_265_p2[32'd44];
        Range2_all_ones_180_reg_11472 <= r_V_199_fu_255_p2[32'd53];
        Range2_all_ones_182_reg_11501 <= r_V_201_fu_257_p2[32'd40];
        Range2_all_ones_183_reg_11530 <= r_V_202_fu_252_p2[32'd53];
        Range2_all_ones_184_reg_11559 <= r_V_203_fu_253_p2[32'd53];
        Range2_all_ones_reg_10793 <= r_V_178_fu_254_p2[32'd42];
        a_V_2_reg_11309 <= {{p_read_int_reg[95:64]}};
        lhs_151_reg_11566 <= lhs_151_fu_7782_p3;
        lhs_152_reg_11572 <= lhs_152_fu_7884_p3;
        lhs_153_reg_11578 <= lhs_153_fu_7986_p3;
        lhs_154_reg_11584 <= lhs_154_fu_8088_p3;
        lhs_155_reg_11590 <= lhs_155_fu_8190_p3;
        lhs_156_reg_11596 <= lhs_156_fu_8292_p3;
        lhs_157_reg_11602 <= lhs_157_fu_8394_p3;
        lhs_158_reg_11608 <= lhs_158_fu_8496_p3;
        lhs_159_reg_11614 <= lhs_159_fu_8598_p3;
        or_ln346_183_reg_11329 <= or_ln346_183_fu_3976_p2;
        or_ln346_183_reg_11329_pp0_iter1_reg <= or_ln346_183_reg_11329;
        overflow_345_reg_11324 <= overflow_345_fu_3946_p2;
        overflow_345_reg_11324_pp0_iter1_reg <= overflow_345_reg_11324;
        p_Result_807_reg_10775 <= r_V_178_fu_254_p2[32'd42];
        p_Result_808_reg_10786 <= p_Val2_807_fu_2783_p2[32'd19];
        p_Result_809_reg_10800 <= r_V_179_fu_262_p2[32'd43];
        p_Result_810_reg_10806 <= r_V_179_fu_262_p2[32'd43];
        p_Result_811_reg_10817 <= p_Val2_810_fu_2847_p2[32'd20];
        p_Result_812_reg_10831 <= r_V_180_fu_251_p2[32'd56];
        p_Result_813_reg_10837 <= r_V_180_fu_251_p2[32'd55];
        p_Result_814_reg_10848 <= p_Val2_813_fu_2907_p2[32'd31];
        p_Result_815_reg_10862 <= r_V_181_fu_256_p2[32'd43];
        p_Result_816_reg_10868 <= r_V_181_fu_256_p2[32'd43];
        p_Result_817_reg_10879 <= p_Val2_816_fu_2971_p2[32'd20];
        p_Result_818_reg_10893 <= r_V_182_fu_264_p2[32'd46];
        p_Result_819_reg_10899 <= r_V_182_fu_264_p2[32'd46];
        p_Result_820_reg_10910 <= p_Val2_819_fu_3035_p2[32'd23];
        p_Result_821_reg_10924 <= r_V_183_fu_240_p2[32'd42];
        p_Result_822_reg_10930 <= r_V_183_fu_240_p2[32'd42];
        p_Result_823_reg_10941 <= p_Val2_822_fu_3099_p2[32'd19];
        p_Result_824_reg_10955 <= r_V_184_fu_249_p2[32'd42];
        p_Result_825_reg_10961 <= r_V_184_fu_249_p2[32'd42];
        p_Result_826_reg_10972 <= p_Val2_825_fu_3163_p2[32'd19];
        p_Result_827_reg_10986 <= r_V_185_fu_259_p2[32'd53];
        p_Result_828_reg_10992 <= r_V_185_fu_259_p2[32'd53];
        p_Result_829_reg_11003 <= p_Val2_828_fu_3227_p2[32'd30];
        p_Result_830_reg_11017 <= r_V_186_fu_246_p2[32'd53];
        p_Result_831_reg_11023 <= r_V_186_fu_246_p2[32'd53];
        p_Result_832_reg_11034 <= p_Val2_831_fu_3291_p2[32'd30];
        p_Result_833_reg_11048 <= r_V_187_fu_266_p2[32'd40];
        p_Result_834_reg_11059 <= r_V_187_fu_266_p2[32'd40];
        p_Result_836_reg_11077 <= r_V_188_fu_261_p2[32'd42];
        p_Result_837_reg_11088 <= r_V_188_fu_261_p2[32'd42];
        p_Result_839_reg_11106 <= r_V_189_fu_242_p2[32'd44];
        p_Result_840_reg_11117 <= r_V_189_fu_242_p2[32'd44];
        p_Result_842_reg_11135 <= r_V_190_fu_260_p2[32'd42];
        p_Result_843_reg_11146 <= r_V_190_fu_260_p2[32'd42];
        p_Result_845_reg_11164 <= r_V_191_fu_263_p2[32'd53];
        p_Result_846_reg_11175 <= r_V_191_fu_263_p2[32'd53];
        p_Result_848_reg_11193 <= r_V_192_fu_250_p2[32'd42];
        p_Result_849_reg_11204 <= r_V_192_fu_250_p2[32'd42];
        p_Result_851_reg_11222 <= r_V_193_fu_244_p2[32'd42];
        p_Result_852_reg_11233 <= r_V_193_fu_244_p2[32'd42];
        p_Result_854_reg_11251 <= r_V_194_fu_243_p2[32'd53];
        p_Result_855_reg_11262 <= r_V_194_fu_243_p2[32'd53];
        p_Result_857_reg_11280 <= r_V_195_fu_248_p2[32'd53];
        p_Result_858_reg_11291 <= r_V_195_fu_248_p2[32'd53];
        p_Result_860_reg_11334 <= r_V_fu_247_p2[32'd42];
        p_Result_861_reg_11345 <= r_V_fu_247_p2[32'd42];
        p_Result_863_reg_11363 <= r_V_196_fu_258_p2[32'd41];
        p_Result_864_reg_11374 <= r_V_196_fu_258_p2[32'd41];
        p_Result_866_reg_11392 <= r_V_197_fu_245_p2[32'd43];
        p_Result_867_reg_11403 <= r_V_197_fu_245_p2[32'd43];
        p_Result_869_reg_11421 <= r_V_198_fu_265_p2[32'd44];
        p_Result_870_reg_11432 <= r_V_198_fu_265_p2[32'd44];
        p_Result_872_reg_11450 <= r_V_199_fu_255_p2[32'd53];
        p_Result_873_reg_11461 <= r_V_199_fu_255_p2[32'd53];
        p_Result_878_reg_11479 <= r_V_201_fu_257_p2[32'd40];
        p_Result_879_reg_11490 <= r_V_201_fu_257_p2[32'd40];
        p_Result_881_reg_11508 <= r_V_202_fu_252_p2[32'd53];
        p_Result_882_reg_11519 <= r_V_202_fu_252_p2[32'd53];
        p_Result_884_reg_11537 <= r_V_203_fu_253_p2[32'd53];
        p_Result_885_reg_11548 <= r_V_203_fu_253_p2[32'd53];
        p_Result_s_reg_10769 <= r_V_178_fu_254_p2[32'd42];
        p_Val2_807_reg_10781 <= p_Val2_807_fu_2783_p2;
        p_Val2_810_reg_10812 <= p_Val2_810_fu_2847_p2;
        p_Val2_813_reg_10843 <= p_Val2_813_fu_2907_p2;
        p_Val2_816_reg_10874 <= p_Val2_816_fu_2971_p2;
        p_Val2_819_reg_10905 <= p_Val2_819_fu_3035_p2;
        p_Val2_822_reg_10936 <= p_Val2_822_fu_3099_p2;
        p_Val2_825_reg_10967 <= p_Val2_825_fu_3163_p2;
        p_Val2_828_reg_10998 <= p_Val2_828_fu_3227_p2;
        p_Val2_831_reg_11029 <= p_Val2_831_fu_3291_p2;
        p_Val2_833_reg_11054 <= {{r_V_187_fu_266_p2[40:24]}};
        p_Val2_836_reg_11083 <= {{r_V_188_fu_261_p2[42:24]}};
        p_Val2_839_reg_11112 <= {{r_V_189_fu_242_p2[44:24]}};
        p_Val2_842_reg_11141 <= {{r_V_190_fu_260_p2[42:24]}};
        p_Val2_845_reg_11170 <= {{r_V_191_fu_263_p2[53:24]}};
        p_Val2_848_reg_11199 <= {{r_V_192_fu_250_p2[42:24]}};
        p_Val2_851_reg_11228 <= {{r_V_193_fu_244_p2[42:24]}};
        p_Val2_854_reg_11257 <= {{r_V_194_fu_243_p2[53:24]}};
        p_Val2_857_reg_11286 <= {{r_V_195_fu_248_p2[53:24]}};
        p_Val2_860_reg_11340 <= {{r_V_fu_247_p2[42:24]}};
        p_Val2_863_reg_11369 <= {{r_V_196_fu_258_p2[41:24]}};
        p_Val2_866_reg_11398 <= {{r_V_197_fu_245_p2[43:24]}};
        p_Val2_869_reg_11427 <= {{r_V_198_fu_265_p2[44:24]}};
        p_Val2_872_reg_11456 <= {{r_V_199_fu_255_p2[53:24]}};
        p_Val2_876_reg_11319 <= p_Val2_876_fu_3844_p2;
        p_Val2_876_reg_11319_pp0_iter1_reg <= p_Val2_876_reg_11319;
        p_Val2_878_reg_11485 <= {{r_V_201_fu_257_p2[40:24]}};
        p_Val2_881_reg_11514 <= {{r_V_202_fu_252_p2[53:24]}};
        p_Val2_884_reg_11543 <= {{r_V_203_fu_253_p2[53:24]}};
        r_V_178_reg_2283 <= r_V_178_fu_254_p2;
        r_V_179_reg_2287 <= r_V_179_fu_262_p2;
        r_V_180_reg_2291 <= r_V_180_fu_251_p2;
        r_V_181_reg_2295 <= r_V_181_fu_256_p2;
        r_V_182_reg_2299 <= r_V_182_fu_264_p2;
        r_V_183_reg_2303 <= r_V_183_fu_240_p2;
        r_V_184_reg_2307 <= r_V_184_fu_249_p2;
        r_V_185_reg_2311 <= r_V_185_fu_259_p2;
        r_V_186_reg_2315 <= r_V_186_fu_246_p2;
        r_V_187_reg_2319 <= r_V_187_fu_266_p2;
        r_V_188_reg_2323 <= r_V_188_fu_261_p2;
        r_V_189_reg_2327 <= r_V_189_fu_242_p2;
        r_V_190_reg_2331 <= r_V_190_fu_260_p2;
        r_V_191_reg_2335 <= r_V_191_fu_263_p2;
        r_V_192_reg_2339 <= r_V_192_fu_250_p2;
        r_V_193_reg_2343 <= r_V_193_fu_244_p2;
        r_V_194_reg_2347 <= r_V_194_fu_243_p2;
        r_V_195_reg_2351 <= r_V_195_fu_248_p2;
        r_V_196_reg_2679 <= r_V_196_fu_258_p2;
        r_V_197_reg_2683 <= r_V_197_fu_245_p2;
        r_V_198_reg_2687 <= r_V_198_fu_265_p2;
        r_V_199_reg_2691 <= r_V_199_fu_255_p2;
        r_V_201_reg_2695 <= r_V_201_fu_257_p2;
        r_V_202_reg_2699 <= r_V_202_fu_252_p2;
        r_V_203_reg_2703 <= r_V_203_fu_253_p2;
        r_V_reg_2675 <= r_V_fu_247_p2;
        tmp_1338_reg_11065 <= r_V_187_fu_266_p2[32'd23];
        tmp_1344_reg_11094 <= r_V_188_fu_261_p2[32'd23];
        tmp_1350_reg_11123 <= r_V_189_fu_242_p2[32'd23];
        tmp_1356_reg_11152 <= r_V_190_fu_260_p2[32'd23];
        tmp_1362_reg_11181 <= r_V_191_fu_263_p2[32'd23];
        tmp_1368_reg_11210 <= r_V_192_fu_250_p2[32'd23];
        tmp_1374_reg_11239 <= r_V_193_fu_244_p2[32'd23];
        tmp_1380_reg_11268 <= r_V_194_fu_243_p2[32'd23];
        tmp_1386_reg_11297 <= r_V_195_fu_248_p2[32'd23];
        tmp_1392_reg_11351 <= r_V_fu_247_p2[32'd23];
        tmp_1398_reg_11380 <= r_V_196_fu_258_p2[32'd23];
        tmp_1404_reg_11409 <= r_V_197_fu_245_p2[32'd23];
        tmp_1410_reg_11438 <= r_V_198_fu_265_p2[32'd23];
        tmp_1416_reg_11467 <= r_V_199_fu_255_p2[32'd23];
        tmp_1428_reg_11496 <= r_V_201_fu_257_p2[32'd23];
        tmp_1434_reg_11525 <= r_V_202_fu_252_p2[32'd23];
        tmp_1440_reg_11554 <= r_V_203_fu_253_p2[32'd23];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= select_ln302_359_fu_9907_p3;
        ap_return_1_int_reg <= select_ln302_361_fu_10007_p3;
        ap_return_2_int_reg <= select_ln302_363_fu_10107_p3;
        ap_return_3_int_reg <= select_ln302_365_fu_10207_p3;
        ap_return_4_int_reg <= select_ln302_367_fu_10307_p3;
        ap_return_5_int_reg <= select_ln302_369_fu_10407_p3;
        ap_return_6_int_reg <= select_ln302_371_fu_10507_p3;
        ap_return_7_int_reg <= select_ln302_373_fu_10607_p3;
        ap_return_8_int_reg <= select_ln302_375_fu_10707_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        p_read_int_reg <= p_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = select_ln302_359_fu_9907_p3;
    end else begin
        ap_return_0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = select_ln302_361_fu_10007_p3;
    end else begin
        ap_return_1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = select_ln302_363_fu_10107_p3;
    end else begin
        ap_return_2 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = select_ln302_365_fu_10207_p3;
    end else begin
        ap_return_3 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = select_ln302_367_fu_10307_p3;
    end else begin
        ap_return_4 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = select_ln302_369_fu_10407_p3;
    end else begin
        ap_return_5 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = select_ln302_371_fu_10507_p3;
    end else begin
        ap_return_6 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = select_ln302_373_fu_10607_p3;
    end else begin
        ap_return_7 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = select_ln302_375_fu_10707_p3;
    end else begin
        ap_return_8 = 'bx;
    end
end

assign Range2_all_ones_181_fu_3870_p3 = r_V_200_fu_3790_p2[32'd38];

assign a_V_1_fu_3313_p4 = {{p_read_int_reg[63:32]}};

assign a_V_2_cast_fu_3736_p4 = {{p_read_int_reg[87:64]}};

assign a_V_2_fu_3726_p4 = {{p_read_int_reg[95:64]}};

assign a_V_fu_2708_p1 = p_read_int_reg[31:0];

assign add_ln823_fu_3818_p2 = (trunc_ln7_fu_3782_p3 + a_V_2_cast_fu_3736_p4);

assign and_ln891_161_fu_4160_p2 = (carry_322_fu_4115_p2 & Range2_all_ones_159_reg_10824);

assign and_ln891_162_fu_4282_p2 = (carry_324_fu_4237_p2 & Range2_all_ones_160_reg_10855);

assign and_ln891_163_fu_4406_p2 = (carry_326_fu_4361_p2 & Range2_all_ones_161_reg_10886);

assign and_ln891_164_fu_4531_p2 = (carry_328_fu_4486_p2 & Range2_all_ones_162_reg_10917);

assign and_ln891_165_fu_4656_p2 = (carry_330_fu_4611_p2 & Range2_all_ones_163_reg_10948);

assign and_ln891_166_fu_4781_p2 = (carry_332_fu_4736_p2 & Range2_all_ones_164_reg_10979);

assign and_ln891_167_fu_4906_p2 = (carry_334_fu_4861_p2 & Range2_all_ones_165_reg_11010);

assign and_ln891_168_fu_5031_p2 = (carry_336_fu_4986_p2 & Range2_all_ones_166_reg_11041);

assign and_ln891_169_fu_5179_p2 = (carry_338_fu_5133_p2 & Range2_all_ones_167_reg_11070);

assign and_ln891_170_fu_5328_p2 = (carry_340_fu_5282_p2 & Range2_all_ones_168_reg_11099);

assign and_ln891_171_fu_5477_p2 = (carry_342_fu_5431_p2 & Range2_all_ones_169_reg_11128);

assign and_ln891_172_fu_5626_p2 = (carry_344_fu_5580_p2 & Range2_all_ones_170_reg_11157);

assign and_ln891_173_fu_5775_p2 = (carry_346_fu_5729_p2 & Range2_all_ones_171_reg_11186);

assign and_ln891_174_fu_5924_p2 = (carry_348_fu_5878_p2 & Range2_all_ones_172_reg_11215);

assign and_ln891_175_fu_6073_p2 = (carry_350_fu_6027_p2 & Range2_all_ones_173_reg_11244);

assign and_ln891_176_fu_6222_p2 = (carry_352_fu_6176_p2 & Range2_all_ones_174_reg_11273);

assign and_ln891_177_fu_6371_p2 = (carry_354_fu_6325_p2 & Range2_all_ones_175_reg_11302);

assign and_ln891_178_fu_8682_p2 = (carry_356_fu_8636_p2 & Range2_all_ones_176_reg_11356);

assign and_ln891_179_fu_8831_p2 = (carry_358_fu_8785_p2 & Range2_all_ones_177_reg_11385);

assign and_ln891_180_fu_8980_p2 = (carry_360_fu_8934_p2 & Range2_all_ones_178_reg_11414);

assign and_ln891_181_fu_9129_p2 = (carry_362_fu_9083_p2 & Range2_all_ones_179_reg_11443);

assign and_ln891_182_fu_9278_p2 = (carry_364_fu_9232_p2 & Range2_all_ones_180_reg_11472);

assign and_ln891_183_fu_3922_p2 = (carry_366_fu_3864_p2 & Range2_all_ones_181_fu_3870_p3);

assign and_ln891_184_fu_9444_p2 = (carry_368_fu_9398_p2 & Range2_all_ones_182_reg_11501);

assign and_ln891_185_fu_9593_p2 = (carry_370_fu_9547_p2 & Range2_all_ones_183_reg_11530);

assign and_ln891_186_fu_9742_p2 = (carry_372_fu_9696_p2 & Range2_all_ones_184_reg_11559);

assign and_ln891_fu_4035_p2 = (carry_320_fu_3990_p2 & Range2_all_ones_reg_10793);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign carry_320_fu_3990_p2 = (xor_ln896_fu_3985_p2 & p_Result_807_reg_10775);

assign carry_322_fu_4115_p2 = (xor_ln896_486_fu_4110_p2 & p_Result_810_reg_10806);

assign carry_324_fu_4237_p2 = (xor_ln896_488_fu_4232_p2 & p_Result_813_reg_10837);

assign carry_326_fu_4361_p2 = (xor_ln896_490_fu_4356_p2 & p_Result_816_reg_10868);

assign carry_328_fu_4486_p2 = (xor_ln896_492_fu_4481_p2 & p_Result_819_reg_10899);

assign carry_330_fu_4611_p2 = (xor_ln896_494_fu_4606_p2 & p_Result_822_reg_10930);

assign carry_332_fu_4736_p2 = (xor_ln896_496_fu_4731_p2 & p_Result_825_reg_10961);

assign carry_334_fu_4861_p2 = (xor_ln896_498_fu_4856_p2 & p_Result_828_reg_10992);

assign carry_336_fu_4986_p2 = (xor_ln896_500_fu_4981_p2 & p_Result_831_reg_11023);

assign carry_338_fu_5133_p2 = (xor_ln896_502_fu_5127_p2 & p_Result_834_reg_11059);

assign carry_340_fu_5282_p2 = (xor_ln896_504_fu_5276_p2 & p_Result_837_reg_11088);

assign carry_342_fu_5431_p2 = (xor_ln896_506_fu_5425_p2 & p_Result_840_reg_11117);

assign carry_344_fu_5580_p2 = (xor_ln896_508_fu_5574_p2 & p_Result_843_reg_11146);

assign carry_346_fu_5729_p2 = (xor_ln896_510_fu_5723_p2 & p_Result_846_reg_11175);

assign carry_348_fu_5878_p2 = (xor_ln896_512_fu_5872_p2 & p_Result_849_reg_11204);

assign carry_350_fu_6027_p2 = (xor_ln896_514_fu_6021_p2 & p_Result_852_reg_11233);

assign carry_352_fu_6176_p2 = (xor_ln896_516_fu_6170_p2 & p_Result_855_reg_11262);

assign carry_354_fu_6325_p2 = (xor_ln896_518_fu_6319_p2 & p_Result_858_reg_11291);

assign carry_356_fu_8636_p2 = (xor_ln896_520_fu_8630_p2 & p_Result_861_reg_11345);

assign carry_358_fu_8785_p2 = (xor_ln896_522_fu_8779_p2 & p_Result_864_reg_11374);

assign carry_360_fu_8934_p2 = (xor_ln896_524_fu_8928_p2 & p_Result_867_reg_11403);

assign carry_362_fu_9083_p2 = (xor_ln896_526_fu_9077_p2 & p_Result_870_reg_11432);

assign carry_364_fu_9232_p2 = (xor_ln896_528_fu_9226_p2 & p_Result_873_reg_11461);

assign carry_366_fu_3864_p2 = (xor_ln896_530_fu_3858_p2 & p_Result_876_fu_3824_p3);

assign carry_368_fu_9398_p2 = (xor_ln896_532_fu_9392_p2 & p_Result_879_reg_11490);

assign carry_370_fu_9547_p2 = (xor_ln896_534_fu_9541_p2 & p_Result_882_reg_11519);

assign carry_372_fu_9696_p2 = (xor_ln896_536_fu_9690_p2 & p_Result_885_reg_11548);

assign deleted_ones_323_fu_4155_p2 = (or_ln890_161_fu_4149_p2 & Range2_all_ones_159_reg_10824);

assign deleted_ones_324_fu_4277_p2 = (or_ln890_162_fu_4271_p2 & Range2_all_ones_160_reg_10855);

assign deleted_ones_325_fu_4401_p2 = (or_ln890_163_fu_4395_p2 & Range2_all_ones_161_reg_10886);

assign deleted_ones_326_fu_4526_p2 = (or_ln890_164_fu_4520_p2 & Range2_all_ones_162_reg_10917);

assign deleted_ones_327_fu_4651_p2 = (or_ln890_165_fu_4645_p2 & Range2_all_ones_163_reg_10948);

assign deleted_ones_328_fu_4776_p2 = (or_ln890_166_fu_4770_p2 & Range2_all_ones_164_reg_10979);

assign deleted_ones_329_fu_4901_p2 = (or_ln890_167_fu_4895_p2 & Range2_all_ones_165_reg_11010);

assign deleted_ones_330_fu_5026_p2 = (or_ln890_168_fu_5020_p2 & Range2_all_ones_166_reg_11041);

assign deleted_ones_331_fu_5174_p2 = (or_ln890_169_fu_5168_p2 & Range2_all_ones_167_reg_11070);

assign deleted_ones_332_fu_5323_p2 = (or_ln890_170_fu_5317_p2 & Range2_all_ones_168_reg_11099);

assign deleted_ones_333_fu_5472_p2 = (or_ln890_171_fu_5466_p2 & Range2_all_ones_169_reg_11128);

assign deleted_ones_334_fu_5621_p2 = (or_ln890_172_fu_5615_p2 & Range2_all_ones_170_reg_11157);

assign deleted_ones_335_fu_5770_p2 = (or_ln890_173_fu_5764_p2 & Range2_all_ones_171_reg_11186);

assign deleted_ones_336_fu_5919_p2 = (or_ln890_174_fu_5913_p2 & Range2_all_ones_172_reg_11215);

assign deleted_ones_337_fu_6068_p2 = (or_ln890_175_fu_6062_p2 & Range2_all_ones_173_reg_11244);

assign deleted_ones_338_fu_6217_p2 = (or_ln890_176_fu_6211_p2 & Range2_all_ones_174_reg_11273);

assign deleted_ones_339_fu_6366_p2 = (or_ln890_177_fu_6360_p2 & Range2_all_ones_175_reg_11302);

assign deleted_ones_340_fu_8677_p2 = (or_ln890_178_fu_8671_p2 & Range2_all_ones_176_reg_11356);

assign deleted_ones_341_fu_8826_p2 = (or_ln890_179_fu_8820_p2 & Range2_all_ones_177_reg_11385);

assign deleted_ones_342_fu_8975_p2 = (or_ln890_180_fu_8969_p2 & Range2_all_ones_178_reg_11414);

assign deleted_ones_343_fu_9124_p2 = (or_ln890_181_fu_9118_p2 & Range2_all_ones_179_reg_11443);

assign deleted_ones_344_fu_9273_p2 = (or_ln890_182_fu_9267_p2 & Range2_all_ones_180_reg_11472);

assign deleted_ones_345_fu_3916_p2 = (or_ln890_183_fu_3910_p2 & Range2_all_ones_181_fu_3870_p3);

assign deleted_ones_346_fu_9439_p2 = (or_ln890_184_fu_9433_p2 & Range2_all_ones_182_reg_11501);

assign deleted_ones_347_fu_9588_p2 = (or_ln890_185_fu_9582_p2 & Range2_all_ones_183_reg_11530);

assign deleted_ones_348_fu_9737_p2 = (or_ln890_186_fu_9731_p2 & Range2_all_ones_184_reg_11559);

assign deleted_ones_fu_4030_p2 = (or_ln890_fu_4024_p2 & Range2_all_ones_reg_10793);

assign deleted_zeros_158_fu_4130_p2 = (or_ln888_161_fu_4125_p2 ^ Range2_all_ones_159_reg_10824);

assign deleted_zeros_159_fu_4252_p2 = (or_ln888_162_fu_4247_p2 ^ Range2_all_ones_160_reg_10855);

assign deleted_zeros_160_fu_4376_p2 = (or_ln888_163_fu_4371_p2 ^ Range2_all_ones_161_reg_10886);

assign deleted_zeros_161_fu_4501_p2 = (or_ln888_164_fu_4496_p2 ^ Range2_all_ones_162_reg_10917);

assign deleted_zeros_162_fu_4626_p2 = (or_ln888_165_fu_4621_p2 ^ Range2_all_ones_163_reg_10948);

assign deleted_zeros_163_fu_4751_p2 = (or_ln888_166_fu_4746_p2 ^ Range2_all_ones_164_reg_10979);

assign deleted_zeros_164_fu_4876_p2 = (or_ln888_167_fu_4871_p2 ^ Range2_all_ones_165_reg_11010);

assign deleted_zeros_165_fu_5001_p2 = (or_ln888_168_fu_4996_p2 ^ Range2_all_ones_166_reg_11041);

assign deleted_zeros_166_fu_5149_p2 = (or_ln888_169_fu_5143_p2 ^ Range2_all_ones_167_reg_11070);

assign deleted_zeros_167_fu_5298_p2 = (or_ln888_170_fu_5292_p2 ^ Range2_all_ones_168_reg_11099);

assign deleted_zeros_168_fu_5447_p2 = (or_ln888_171_fu_5441_p2 ^ Range2_all_ones_169_reg_11128);

assign deleted_zeros_169_fu_5596_p2 = (or_ln888_172_fu_5590_p2 ^ Range2_all_ones_170_reg_11157);

assign deleted_zeros_170_fu_5745_p2 = (or_ln888_173_fu_5739_p2 ^ Range2_all_ones_171_reg_11186);

assign deleted_zeros_171_fu_5894_p2 = (or_ln888_174_fu_5888_p2 ^ Range2_all_ones_172_reg_11215);

assign deleted_zeros_172_fu_6043_p2 = (or_ln888_175_fu_6037_p2 ^ Range2_all_ones_173_reg_11244);

assign deleted_zeros_173_fu_6192_p2 = (or_ln888_176_fu_6186_p2 ^ Range2_all_ones_174_reg_11273);

assign deleted_zeros_174_fu_6341_p2 = (or_ln888_177_fu_6335_p2 ^ Range2_all_ones_175_reg_11302);

assign deleted_zeros_175_fu_8652_p2 = (or_ln888_178_fu_8646_p2 ^ Range2_all_ones_176_reg_11356);

assign deleted_zeros_176_fu_8801_p2 = (or_ln888_179_fu_8795_p2 ^ Range2_all_ones_177_reg_11385);

assign deleted_zeros_177_fu_8950_p2 = (or_ln888_180_fu_8944_p2 ^ Range2_all_ones_178_reg_11414);

assign deleted_zeros_178_fu_9099_p2 = (or_ln888_181_fu_9093_p2 ^ Range2_all_ones_179_reg_11443);

assign deleted_zeros_179_fu_9248_p2 = (or_ln888_182_fu_9242_p2 ^ Range2_all_ones_180_reg_11472);

assign deleted_zeros_180_fu_3890_p2 = (or_ln888_183_fu_3884_p2 ^ Range2_all_ones_181_fu_3870_p3);

assign deleted_zeros_181_fu_9414_p2 = (or_ln888_184_fu_9408_p2 ^ Range2_all_ones_182_reg_11501);

assign deleted_zeros_182_fu_9563_p2 = (or_ln888_185_fu_9557_p2 ^ Range2_all_ones_183_reg_11530);

assign deleted_zeros_183_fu_9712_p2 = (or_ln888_186_fu_9706_p2 ^ Range2_all_ones_184_reg_11559);

assign deleted_zeros_fu_4005_p2 = (or_ln888_fu_4000_p2 ^ Range2_all_ones_reg_10793);

assign lhs_143_fu_6994_p3 = ((or_ln302_161_fu_6972_p2[0:0] == 1'b1) ? select_ln302_324_fu_6978_p3 : select_ln350_161_fu_6986_p3);

assign lhs_144_fu_7092_p3 = ((or_ln302_162_fu_7070_p2[0:0] == 1'b1) ? select_ln302_326_fu_7076_p3 : select_ln350_162_fu_7084_p3);

assign lhs_145_fu_7190_p3 = ((or_ln302_163_fu_7168_p2[0:0] == 1'b1) ? select_ln302_328_fu_7174_p3 : select_ln350_163_fu_7182_p3);

assign lhs_146_fu_7288_p3 = ((or_ln302_164_fu_7266_p2[0:0] == 1'b1) ? select_ln302_330_fu_7272_p3 : select_ln350_164_fu_7280_p3);

assign lhs_147_fu_7386_p3 = ((or_ln302_165_fu_7364_p2[0:0] == 1'b1) ? select_ln302_332_fu_7370_p3 : select_ln350_165_fu_7378_p3);

assign lhs_148_fu_7484_p3 = ((or_ln302_166_fu_7462_p2[0:0] == 1'b1) ? select_ln302_334_fu_7468_p3 : select_ln350_166_fu_7476_p3);

assign lhs_149_fu_7582_p3 = ((or_ln302_167_fu_7560_p2[0:0] == 1'b1) ? select_ln302_336_fu_7566_p3 : select_ln350_167_fu_7574_p3);

assign lhs_150_fu_7680_p3 = ((or_ln302_168_fu_7658_p2[0:0] == 1'b1) ? select_ln302_338_fu_7664_p3 : select_ln350_168_fu_7672_p3);

assign lhs_151_fu_7782_p3 = ((or_ln302_169_fu_7760_p2[0:0] == 1'b1) ? select_ln302_340_fu_7766_p3 : select_ln350_169_fu_7774_p3);

assign lhs_152_fu_7884_p3 = ((or_ln302_170_fu_7862_p2[0:0] == 1'b1) ? select_ln302_342_fu_7868_p3 : select_ln350_170_fu_7876_p3);

assign lhs_153_fu_7986_p3 = ((or_ln302_171_fu_7964_p2[0:0] == 1'b1) ? select_ln302_344_fu_7970_p3 : select_ln350_171_fu_7978_p3);

assign lhs_154_fu_8088_p3 = ((or_ln302_172_fu_8066_p2[0:0] == 1'b1) ? select_ln302_346_fu_8072_p3 : select_ln350_172_fu_8080_p3);

assign lhs_155_fu_8190_p3 = ((or_ln302_173_fu_8168_p2[0:0] == 1'b1) ? select_ln302_348_fu_8174_p3 : select_ln350_173_fu_8182_p3);

assign lhs_156_fu_8292_p3 = ((or_ln302_174_fu_8270_p2[0:0] == 1'b1) ? select_ln302_350_fu_8276_p3 : select_ln350_174_fu_8284_p3);

assign lhs_157_fu_8394_p3 = ((or_ln302_175_fu_8372_p2[0:0] == 1'b1) ? select_ln302_352_fu_8378_p3 : select_ln350_175_fu_8386_p3);

assign lhs_158_fu_8496_p3 = ((or_ln302_176_fu_8474_p2[0:0] == 1'b1) ? select_ln302_354_fu_8480_p3 : select_ln350_176_fu_8488_p3);

assign lhs_159_fu_8598_p3 = ((or_ln302_177_fu_8576_p2[0:0] == 1'b1) ? select_ln302_356_fu_8582_p3 : select_ln350_177_fu_8590_p3);

assign lhs_fu_6896_p3 = ((or_ln302_fu_6874_p2[0:0] == 1'b1) ? select_ln302_fu_6880_p3 : select_ln350_fu_6888_p3);

assign or_ln302_161_fu_6972_p2 = (xor_ln302_325_fu_6966_p2 | overflow_350_fu_6942_p2);

assign or_ln302_162_fu_7070_p2 = (xor_ln302_327_fu_7064_p2 | overflow_351_fu_7040_p2);

assign or_ln302_163_fu_7168_p2 = (xor_ln302_329_fu_7162_p2 | overflow_352_fu_7138_p2);

assign or_ln302_164_fu_7266_p2 = (xor_ln302_331_fu_7260_p2 | overflow_353_fu_7236_p2);

assign or_ln302_165_fu_7364_p2 = (xor_ln302_333_fu_7358_p2 | overflow_354_fu_7334_p2);

assign or_ln302_166_fu_7462_p2 = (xor_ln302_335_fu_7456_p2 | overflow_355_fu_7432_p2);

assign or_ln302_167_fu_7560_p2 = (xor_ln302_337_fu_7554_p2 | overflow_356_fu_7530_p2);

assign or_ln302_168_fu_7658_p2 = (xor_ln302_339_fu_7652_p2 | overflow_357_fu_7628_p2);

assign or_ln302_169_fu_7760_p2 = (xor_ln302_341_fu_7754_p2 | overflow_358_fu_7730_p2);

assign or_ln302_170_fu_7862_p2 = (xor_ln302_343_fu_7856_p2 | overflow_359_fu_7832_p2);

assign or_ln302_171_fu_7964_p2 = (xor_ln302_345_fu_7958_p2 | overflow_360_fu_7934_p2);

assign or_ln302_172_fu_8066_p2 = (xor_ln302_347_fu_8060_p2 | overflow_361_fu_8036_p2);

assign or_ln302_173_fu_8168_p2 = (xor_ln302_349_fu_8162_p2 | overflow_362_fu_8138_p2);

assign or_ln302_174_fu_8270_p2 = (xor_ln302_351_fu_8264_p2 | overflow_363_fu_8240_p2);

assign or_ln302_175_fu_8372_p2 = (xor_ln302_353_fu_8366_p2 | overflow_364_fu_8342_p2);

assign or_ln302_176_fu_8474_p2 = (xor_ln302_355_fu_8468_p2 | overflow_365_fu_8444_p2);

assign or_ln302_177_fu_8576_p2 = (xor_ln302_357_fu_8570_p2 | overflow_366_fu_8546_p2);

assign or_ln302_178_fu_9885_p2 = (xor_ln302_359_fu_9879_p2 | overflow_367_fu_9855_p2);

assign or_ln302_179_fu_9985_p2 = (xor_ln302_361_fu_9979_p2 | overflow_368_fu_9955_p2);

assign or_ln302_180_fu_10085_p2 = (xor_ln302_363_fu_10079_p2 | overflow_369_fu_10055_p2);

assign or_ln302_181_fu_10185_p2 = (xor_ln302_365_fu_10179_p2 | overflow_370_fu_10155_p2);

assign or_ln302_182_fu_10285_p2 = (xor_ln302_367_fu_10279_p2 | overflow_371_fu_10255_p2);

assign or_ln302_183_fu_10385_p2 = (xor_ln302_369_fu_10379_p2 | overflow_372_fu_10355_p2);

assign or_ln302_184_fu_10485_p2 = (xor_ln302_371_fu_10479_p2 | overflow_373_fu_10455_p2);

assign or_ln302_185_fu_10585_p2 = (xor_ln302_373_fu_10579_p2 | overflow_374_fu_10555_p2);

assign or_ln302_186_fu_10685_p2 = (xor_ln302_375_fu_10679_p2 | overflow_375_fu_10655_p2);

assign or_ln302_fu_6874_p2 = (xor_ln302_323_fu_6868_p2 | overflow_349_fu_6844_p2);

assign or_ln346_161_fu_4218_p2 = (underflow_323_fu_4205_p2 | overflow_323_fu_4181_p2);

assign or_ln346_162_fu_4340_p2 = (underflow_324_fu_4327_p2 | overflow_324_fu_4303_p2);

assign or_ln346_163_fu_4464_p2 = (underflow_325_fu_4451_p2 | overflow_325_fu_4427_p2);

assign or_ln346_164_fu_4589_p2 = (underflow_326_fu_4576_p2 | overflow_326_fu_4552_p2);

assign or_ln346_165_fu_4714_p2 = (underflow_327_fu_4701_p2 | overflow_327_fu_4677_p2);

assign or_ln346_166_fu_4839_p2 = (underflow_328_fu_4826_p2 | overflow_328_fu_4802_p2);

assign or_ln346_167_fu_4964_p2 = (underflow_329_fu_4951_p2 | overflow_329_fu_4927_p2);

assign or_ln346_168_fu_5089_p2 = (underflow_330_fu_5076_p2 | overflow_330_fu_5052_p2);

assign or_ln346_169_fu_5238_p2 = (underflow_331_fu_5225_p2 | overflow_331_fu_5201_p2);

assign or_ln346_170_fu_5387_p2 = (underflow_332_fu_5374_p2 | overflow_332_fu_5350_p2);

assign or_ln346_171_fu_5536_p2 = (underflow_333_fu_5523_p2 | overflow_333_fu_5499_p2);

assign or_ln346_172_fu_5685_p2 = (underflow_334_fu_5672_p2 | overflow_334_fu_5648_p2);

assign or_ln346_173_fu_5834_p2 = (underflow_335_fu_5821_p2 | overflow_335_fu_5797_p2);

assign or_ln346_174_fu_5983_p2 = (underflow_336_fu_5970_p2 | overflow_336_fu_5946_p2);

assign or_ln346_175_fu_6132_p2 = (underflow_337_fu_6119_p2 | overflow_337_fu_6095_p2);

assign or_ln346_176_fu_6281_p2 = (underflow_338_fu_6268_p2 | overflow_338_fu_6244_p2);

assign or_ln346_177_fu_6430_p2 = (underflow_339_fu_6417_p2 | overflow_339_fu_6393_p2);

assign or_ln346_178_fu_8741_p2 = (underflow_340_fu_8728_p2 | overflow_340_fu_8704_p2);

assign or_ln346_179_fu_8890_p2 = (underflow_341_fu_8877_p2 | overflow_341_fu_8853_p2);

assign or_ln346_180_fu_9039_p2 = (underflow_342_fu_9026_p2 | overflow_342_fu_9002_p2);

assign or_ln346_181_fu_9188_p2 = (underflow_343_fu_9175_p2 | overflow_343_fu_9151_p2);

assign or_ln346_182_fu_9337_p2 = (underflow_344_fu_9324_p2 | overflow_344_fu_9300_p2);

assign or_ln346_183_fu_3976_p2 = (underflow_345_fu_3970_p2 | overflow_345_fu_3946_p2);

assign or_ln346_184_fu_9503_p2 = (underflow_346_fu_9490_p2 | overflow_346_fu_9466_p2);

assign or_ln346_185_fu_9652_p2 = (underflow_347_fu_9639_p2 | overflow_347_fu_9615_p2);

assign or_ln346_186_fu_9801_p2 = (underflow_348_fu_9788_p2 | overflow_348_fu_9764_p2);

assign or_ln346_fu_4093_p2 = (underflow_fu_4080_p2 | overflow_fu_4056_p2);

assign or_ln888_161_fu_4125_p2 = (xor_ln888_321_fu_4120_p2 | p_Result_811_reg_10817);

assign or_ln888_162_fu_4247_p2 = (xor_ln888_323_fu_4242_p2 | p_Result_814_reg_10848);

assign or_ln888_163_fu_4371_p2 = (xor_ln888_325_fu_4366_p2 | p_Result_817_reg_10879);

assign or_ln888_164_fu_4496_p2 = (xor_ln888_327_fu_4491_p2 | p_Result_820_reg_10910);

assign or_ln888_165_fu_4621_p2 = (xor_ln888_329_fu_4616_p2 | p_Result_823_reg_10941);

assign or_ln888_166_fu_4746_p2 = (xor_ln888_331_fu_4741_p2 | p_Result_826_reg_10972);

assign or_ln888_167_fu_4871_p2 = (xor_ln888_333_fu_4866_p2 | p_Result_829_reg_11003);

assign or_ln888_168_fu_4996_p2 = (xor_ln888_335_fu_4991_p2 | p_Result_832_reg_11034);

assign or_ln888_169_fu_5143_p2 = (xor_ln888_337_fu_5138_p2 | p_Result_835_fu_5119_p3);

assign or_ln888_170_fu_5292_p2 = (xor_ln888_339_fu_5287_p2 | p_Result_838_fu_5268_p3);

assign or_ln888_171_fu_5441_p2 = (xor_ln888_341_fu_5436_p2 | p_Result_841_fu_5417_p3);

assign or_ln888_172_fu_5590_p2 = (xor_ln888_343_fu_5585_p2 | p_Result_844_fu_5566_p3);

assign or_ln888_173_fu_5739_p2 = (xor_ln888_345_fu_5734_p2 | p_Result_847_fu_5715_p3);

assign or_ln888_174_fu_5888_p2 = (xor_ln888_347_fu_5883_p2 | p_Result_850_fu_5864_p3);

assign or_ln888_175_fu_6037_p2 = (xor_ln888_349_fu_6032_p2 | p_Result_853_fu_6013_p3);

assign or_ln888_176_fu_6186_p2 = (xor_ln888_351_fu_6181_p2 | p_Result_856_fu_6162_p3);

assign or_ln888_177_fu_6335_p2 = (xor_ln888_353_fu_6330_p2 | p_Result_859_fu_6311_p3);

assign or_ln888_178_fu_8646_p2 = (xor_ln888_355_fu_8641_p2 | p_Result_862_fu_8622_p3);

assign or_ln888_179_fu_8795_p2 = (xor_ln888_357_fu_8790_p2 | p_Result_865_fu_8771_p3);

assign or_ln888_180_fu_8944_p2 = (xor_ln888_359_fu_8939_p2 | p_Result_868_fu_8920_p3);

assign or_ln888_181_fu_9093_p2 = (xor_ln888_361_fu_9088_p2 | p_Result_871_fu_9069_p3);

assign or_ln888_182_fu_9242_p2 = (xor_ln888_363_fu_9237_p2 | p_Result_874_fu_9218_p3);

assign or_ln888_183_fu_3884_p2 = (xor_ln888_365_fu_3878_p2 | p_Result_877_fu_3850_p3);

assign or_ln888_184_fu_9408_p2 = (xor_ln888_367_fu_9403_p2 | p_Result_880_fu_9384_p3);

assign or_ln888_185_fu_9557_p2 = (xor_ln888_369_fu_9552_p2 | p_Result_883_fu_9533_p3);

assign or_ln888_186_fu_9706_p2 = (xor_ln888_371_fu_9701_p2 | p_Result_886_fu_9682_p3);

assign or_ln888_fu_4000_p2 = (xor_ln888_fu_3995_p2 | p_Result_808_reg_10786);

assign or_ln890_161_fu_4149_p2 = (xor_ln890_159_fu_4143_p2 | or_ln888_161_fu_4125_p2);

assign or_ln890_162_fu_4271_p2 = (xor_ln890_160_fu_4265_p2 | or_ln888_162_fu_4247_p2);

assign or_ln890_163_fu_4395_p2 = (xor_ln890_161_fu_4389_p2 | or_ln888_163_fu_4371_p2);

assign or_ln890_164_fu_4520_p2 = (xor_ln890_162_fu_4514_p2 | or_ln888_164_fu_4496_p2);

assign or_ln890_165_fu_4645_p2 = (xor_ln890_163_fu_4639_p2 | or_ln888_165_fu_4621_p2);

assign or_ln890_166_fu_4770_p2 = (xor_ln890_164_fu_4764_p2 | or_ln888_166_fu_4746_p2);

assign or_ln890_167_fu_4895_p2 = (xor_ln890_165_fu_4889_p2 | or_ln888_167_fu_4871_p2);

assign or_ln890_168_fu_5020_p2 = (xor_ln890_166_fu_5014_p2 | or_ln888_168_fu_4996_p2);

assign or_ln890_169_fu_5168_p2 = (xor_ln890_167_fu_5162_p2 | or_ln888_169_fu_5143_p2);

assign or_ln890_170_fu_5317_p2 = (xor_ln890_168_fu_5311_p2 | or_ln888_170_fu_5292_p2);

assign or_ln890_171_fu_5466_p2 = (xor_ln890_169_fu_5460_p2 | or_ln888_171_fu_5441_p2);

assign or_ln890_172_fu_5615_p2 = (xor_ln890_170_fu_5609_p2 | or_ln888_172_fu_5590_p2);

assign or_ln890_173_fu_5764_p2 = (xor_ln890_171_fu_5758_p2 | or_ln888_173_fu_5739_p2);

assign or_ln890_174_fu_5913_p2 = (xor_ln890_172_fu_5907_p2 | or_ln888_174_fu_5888_p2);

assign or_ln890_175_fu_6062_p2 = (xor_ln890_173_fu_6056_p2 | or_ln888_175_fu_6037_p2);

assign or_ln890_176_fu_6211_p2 = (xor_ln890_174_fu_6205_p2 | or_ln888_176_fu_6186_p2);

assign or_ln890_177_fu_6360_p2 = (xor_ln890_175_fu_6354_p2 | or_ln888_177_fu_6335_p2);

assign or_ln890_178_fu_8671_p2 = (xor_ln890_176_fu_8665_p2 | or_ln888_178_fu_8646_p2);

assign or_ln890_179_fu_8820_p2 = (xor_ln890_177_fu_8814_p2 | or_ln888_179_fu_8795_p2);

assign or_ln890_180_fu_8969_p2 = (xor_ln890_178_fu_8963_p2 | or_ln888_180_fu_8944_p2);

assign or_ln890_181_fu_9118_p2 = (xor_ln890_179_fu_9112_p2 | or_ln888_181_fu_9093_p2);

assign or_ln890_182_fu_9267_p2 = (xor_ln890_180_fu_9261_p2 | or_ln888_182_fu_9242_p2);

assign or_ln890_183_fu_3910_p2 = (xor_ln890_181_fu_3904_p2 | or_ln888_183_fu_3884_p2);

assign or_ln890_184_fu_9433_p2 = (xor_ln890_182_fu_9427_p2 | or_ln888_184_fu_9408_p2);

assign or_ln890_185_fu_9582_p2 = (xor_ln890_183_fu_9576_p2 | or_ln888_185_fu_9557_p2);

assign or_ln890_186_fu_9731_p2 = (xor_ln890_184_fu_9725_p2 | or_ln888_186_fu_9706_p2);

assign or_ln890_fu_4024_p2 = (xor_ln890_fu_4018_p2 | or_ln888_fu_4000_p2);

assign or_ln895_161_fu_4171_p2 = (xor_ln895_486_fu_4165_p2 | p_Result_811_reg_10817);

assign or_ln895_162_fu_4293_p2 = (xor_ln895_488_fu_4287_p2 | p_Result_814_reg_10848);

assign or_ln895_163_fu_4417_p2 = (xor_ln895_490_fu_4411_p2 | p_Result_817_reg_10879);

assign or_ln895_164_fu_4542_p2 = (xor_ln895_492_fu_4536_p2 | p_Result_820_reg_10910);

assign or_ln895_165_fu_4667_p2 = (xor_ln895_494_fu_4661_p2 | p_Result_823_reg_10941);

assign or_ln895_166_fu_4792_p2 = (xor_ln895_496_fu_4786_p2 | p_Result_826_reg_10972);

assign or_ln895_167_fu_4917_p2 = (xor_ln895_498_fu_4911_p2 | p_Result_829_reg_11003);

assign or_ln895_168_fu_5042_p2 = (xor_ln895_500_fu_5036_p2 | p_Result_832_reg_11034);

assign or_ln895_169_fu_5190_p2 = (xor_ln895_502_fu_5184_p2 | p_Result_835_fu_5119_p3);

assign or_ln895_170_fu_5339_p2 = (xor_ln895_504_fu_5333_p2 | p_Result_838_fu_5268_p3);

assign or_ln895_171_fu_5488_p2 = (xor_ln895_506_fu_5482_p2 | p_Result_841_fu_5417_p3);

assign or_ln895_172_fu_5637_p2 = (xor_ln895_508_fu_5631_p2 | p_Result_844_fu_5566_p3);

assign or_ln895_173_fu_5786_p2 = (xor_ln895_510_fu_5780_p2 | p_Result_847_fu_5715_p3);

assign or_ln895_174_fu_5935_p2 = (xor_ln895_512_fu_5929_p2 | p_Result_850_fu_5864_p3);

assign or_ln895_175_fu_6084_p2 = (xor_ln895_514_fu_6078_p2 | p_Result_853_fu_6013_p3);

assign or_ln895_176_fu_6233_p2 = (xor_ln895_516_fu_6227_p2 | p_Result_856_fu_6162_p3);

assign or_ln895_177_fu_6382_p2 = (xor_ln895_518_fu_6376_p2 | p_Result_859_fu_6311_p3);

assign or_ln895_178_fu_8693_p2 = (xor_ln895_520_fu_8687_p2 | p_Result_862_fu_8622_p3);

assign or_ln895_179_fu_8842_p2 = (xor_ln895_522_fu_8836_p2 | p_Result_865_fu_8771_p3);

assign or_ln895_180_fu_8991_p2 = (xor_ln895_524_fu_8985_p2 | p_Result_868_fu_8920_p3);

assign or_ln895_181_fu_9140_p2 = (xor_ln895_526_fu_9134_p2 | p_Result_871_fu_9069_p3);

assign or_ln895_182_fu_9289_p2 = (xor_ln895_528_fu_9283_p2 | p_Result_874_fu_9218_p3);

assign or_ln895_183_fu_3934_p2 = (xor_ln895_530_fu_3928_p2 | p_Result_877_fu_3850_p3);

assign or_ln895_184_fu_9455_p2 = (xor_ln895_532_fu_9449_p2 | p_Result_880_fu_9384_p3);

assign or_ln895_185_fu_9604_p2 = (xor_ln895_534_fu_9598_p2 | p_Result_883_fu_9533_p3);

assign or_ln895_186_fu_9753_p2 = (xor_ln895_536_fu_9747_p2 | p_Result_886_fu_9682_p3);

assign or_ln895_fu_4046_p2 = (xor_ln895_fu_4040_p2 | p_Result_808_reg_10786);

assign or_ln896_161_fu_4193_p2 = (xor_ln896_487_fu_4187_p2 | xor_ln896_486_fu_4110_p2);

assign or_ln896_162_fu_4315_p2 = (xor_ln896_489_fu_4309_p2 | xor_ln896_488_fu_4232_p2);

assign or_ln896_163_fu_4439_p2 = (xor_ln896_491_fu_4433_p2 | xor_ln896_490_fu_4356_p2);

assign or_ln896_164_fu_4564_p2 = (xor_ln896_493_fu_4558_p2 | xor_ln896_492_fu_4481_p2);

assign or_ln896_165_fu_4689_p2 = (xor_ln896_495_fu_4683_p2 | xor_ln896_494_fu_4606_p2);

assign or_ln896_166_fu_4814_p2 = (xor_ln896_497_fu_4808_p2 | xor_ln896_496_fu_4731_p2);

assign or_ln896_167_fu_4939_p2 = (xor_ln896_499_fu_4933_p2 | xor_ln896_498_fu_4856_p2);

assign or_ln896_168_fu_5064_p2 = (xor_ln896_501_fu_5058_p2 | xor_ln896_500_fu_4981_p2);

assign or_ln896_169_fu_5213_p2 = (xor_ln896_503_fu_5207_p2 | xor_ln896_502_fu_5127_p2);

assign or_ln896_170_fu_5362_p2 = (xor_ln896_505_fu_5356_p2 | xor_ln896_504_fu_5276_p2);

assign or_ln896_171_fu_5511_p2 = (xor_ln896_507_fu_5505_p2 | xor_ln896_506_fu_5425_p2);

assign or_ln896_172_fu_5660_p2 = (xor_ln896_509_fu_5654_p2 | xor_ln896_508_fu_5574_p2);

assign or_ln896_173_fu_5809_p2 = (xor_ln896_511_fu_5803_p2 | xor_ln896_510_fu_5723_p2);

assign or_ln896_174_fu_5958_p2 = (xor_ln896_513_fu_5952_p2 | xor_ln896_512_fu_5872_p2);

assign or_ln896_175_fu_6107_p2 = (xor_ln896_515_fu_6101_p2 | xor_ln896_514_fu_6021_p2);

assign or_ln896_176_fu_6256_p2 = (xor_ln896_517_fu_6250_p2 | xor_ln896_516_fu_6170_p2);

assign or_ln896_177_fu_6405_p2 = (xor_ln896_519_fu_6399_p2 | xor_ln896_518_fu_6319_p2);

assign or_ln896_178_fu_8716_p2 = (xor_ln896_521_fu_8710_p2 | xor_ln896_520_fu_8630_p2);

assign or_ln896_179_fu_8865_p2 = (xor_ln896_523_fu_8859_p2 | xor_ln896_522_fu_8779_p2);

assign or_ln896_180_fu_9014_p2 = (xor_ln896_525_fu_9008_p2 | xor_ln896_524_fu_8928_p2);

assign or_ln896_181_fu_9163_p2 = (xor_ln896_527_fu_9157_p2 | xor_ln896_526_fu_9077_p2);

assign or_ln896_182_fu_9312_p2 = (xor_ln896_529_fu_9306_p2 | xor_ln896_528_fu_9226_p2);

assign or_ln896_183_fu_3958_p2 = (xor_ln896_531_fu_3952_p2 | xor_ln896_530_fu_3858_p2);

assign or_ln896_184_fu_9478_p2 = (xor_ln896_533_fu_9472_p2 | xor_ln896_532_fu_9392_p2);

assign or_ln896_185_fu_9627_p2 = (xor_ln896_535_fu_9621_p2 | xor_ln896_534_fu_9541_p2);

assign or_ln896_186_fu_9776_p2 = (xor_ln896_537_fu_9770_p2 | xor_ln896_536_fu_9690_p2);

assign or_ln896_fu_4068_p2 = (xor_ln896_fu_3985_p2 | xor_ln896_485_fu_4062_p2);

assign overflow_323_fu_4181_p2 = (xor_ln895_487_fu_4176_p2 & or_ln895_161_fu_4171_p2);

assign overflow_324_fu_4303_p2 = (xor_ln895_489_fu_4298_p2 & or_ln895_162_fu_4293_p2);

assign overflow_325_fu_4427_p2 = (xor_ln895_491_fu_4422_p2 & or_ln895_163_fu_4417_p2);

assign overflow_326_fu_4552_p2 = (xor_ln895_493_fu_4547_p2 & or_ln895_164_fu_4542_p2);

assign overflow_327_fu_4677_p2 = (xor_ln895_495_fu_4672_p2 & or_ln895_165_fu_4667_p2);

assign overflow_328_fu_4802_p2 = (xor_ln895_497_fu_4797_p2 & or_ln895_166_fu_4792_p2);

assign overflow_329_fu_4927_p2 = (xor_ln895_499_fu_4922_p2 & or_ln895_167_fu_4917_p2);

assign overflow_330_fu_5052_p2 = (xor_ln895_501_fu_5047_p2 & or_ln895_168_fu_5042_p2);

assign overflow_331_fu_5201_p2 = (xor_ln895_503_fu_5196_p2 & or_ln895_169_fu_5190_p2);

assign overflow_332_fu_5350_p2 = (xor_ln895_505_fu_5345_p2 & or_ln895_170_fu_5339_p2);

assign overflow_333_fu_5499_p2 = (xor_ln895_507_fu_5494_p2 & or_ln895_171_fu_5488_p2);

assign overflow_334_fu_5648_p2 = (xor_ln895_509_fu_5643_p2 & or_ln895_172_fu_5637_p2);

assign overflow_335_fu_5797_p2 = (xor_ln895_511_fu_5792_p2 & or_ln895_173_fu_5786_p2);

assign overflow_336_fu_5946_p2 = (xor_ln895_513_fu_5941_p2 & or_ln895_174_fu_5935_p2);

assign overflow_337_fu_6095_p2 = (xor_ln895_515_fu_6090_p2 & or_ln895_175_fu_6084_p2);

assign overflow_338_fu_6244_p2 = (xor_ln895_517_fu_6239_p2 & or_ln895_176_fu_6233_p2);

assign overflow_339_fu_6393_p2 = (xor_ln895_519_fu_6388_p2 & or_ln895_177_fu_6382_p2);

assign overflow_340_fu_8704_p2 = (xor_ln895_521_fu_8699_p2 & or_ln895_178_fu_8693_p2);

assign overflow_341_fu_8853_p2 = (xor_ln895_523_fu_8848_p2 & or_ln895_179_fu_8842_p2);

assign overflow_342_fu_9002_p2 = (xor_ln895_525_fu_8997_p2 & or_ln895_180_fu_8991_p2);

assign overflow_343_fu_9151_p2 = (xor_ln895_527_fu_9146_p2 & or_ln895_181_fu_9140_p2);

assign overflow_344_fu_9300_p2 = (xor_ln895_529_fu_9295_p2 & or_ln895_182_fu_9289_p2);

assign overflow_345_fu_3946_p2 = (xor_ln895_531_fu_3940_p2 & or_ln895_183_fu_3934_p2);

assign overflow_346_fu_9466_p2 = (xor_ln895_533_fu_9461_p2 & or_ln895_184_fu_9455_p2);

assign overflow_347_fu_9615_p2 = (xor_ln895_535_fu_9610_p2 & or_ln895_185_fu_9604_p2);

assign overflow_348_fu_9764_p2 = (xor_ln895_537_fu_9759_p2 & or_ln895_186_fu_9753_p2);

assign overflow_349_fu_6844_p2 = (xor_ln895_538_fu_6838_p2 & p_Result_888_fu_6830_p3);

assign overflow_350_fu_6942_p2 = (xor_ln895_539_fu_6936_p2 & p_Result_890_fu_6928_p3);

assign overflow_351_fu_7040_p2 = (xor_ln895_540_fu_7034_p2 & p_Result_892_fu_7026_p3);

assign overflow_352_fu_7138_p2 = (xor_ln895_541_fu_7132_p2 & p_Result_894_fu_7124_p3);

assign overflow_353_fu_7236_p2 = (xor_ln895_542_fu_7230_p2 & p_Result_896_fu_7222_p3);

assign overflow_354_fu_7334_p2 = (xor_ln895_543_fu_7328_p2 & p_Result_898_fu_7320_p3);

assign overflow_355_fu_7432_p2 = (xor_ln895_544_fu_7426_p2 & p_Result_900_fu_7418_p3);

assign overflow_356_fu_7530_p2 = (xor_ln895_545_fu_7524_p2 & p_Result_902_fu_7516_p3);

assign overflow_357_fu_7628_p2 = (xor_ln895_546_fu_7622_p2 & p_Result_904_fu_7614_p3);

assign overflow_358_fu_7730_p2 = (xor_ln895_547_fu_7724_p2 & p_Result_906_fu_7716_p3);

assign overflow_359_fu_7832_p2 = (xor_ln895_548_fu_7826_p2 & p_Result_908_fu_7818_p3);

assign overflow_360_fu_7934_p2 = (xor_ln895_549_fu_7928_p2 & p_Result_910_fu_7920_p3);

assign overflow_361_fu_8036_p2 = (xor_ln895_550_fu_8030_p2 & p_Result_912_fu_8022_p3);

assign overflow_362_fu_8138_p2 = (xor_ln895_551_fu_8132_p2 & p_Result_914_fu_8124_p3);

assign overflow_363_fu_8240_p2 = (xor_ln895_552_fu_8234_p2 & p_Result_916_fu_8226_p3);

assign overflow_364_fu_8342_p2 = (xor_ln895_553_fu_8336_p2 & p_Result_918_fu_8328_p3);

assign overflow_365_fu_8444_p2 = (xor_ln895_554_fu_8438_p2 & p_Result_920_fu_8430_p3);

assign overflow_366_fu_8546_p2 = (xor_ln895_555_fu_8540_p2 & p_Result_922_fu_8532_p3);

assign overflow_367_fu_9855_p2 = (xor_ln895_556_fu_9849_p2 & p_Result_924_fu_9841_p3);

assign overflow_368_fu_9955_p2 = (xor_ln895_557_fu_9949_p2 & p_Result_926_fu_9941_p3);

assign overflow_369_fu_10055_p2 = (xor_ln895_558_fu_10049_p2 & p_Result_928_fu_10041_p3);

assign overflow_370_fu_10155_p2 = (xor_ln895_559_fu_10149_p2 & p_Result_930_fu_10141_p3);

assign overflow_371_fu_10255_p2 = (xor_ln895_560_fu_10249_p2 & p_Result_932_fu_10241_p3);

assign overflow_372_fu_10355_p2 = (xor_ln895_561_fu_10349_p2 & p_Result_934_fu_10341_p3);

assign overflow_373_fu_10455_p2 = (xor_ln895_562_fu_10449_p2 & p_Result_936_fu_10441_p3);

assign overflow_374_fu_10555_p2 = (xor_ln895_563_fu_10549_p2 & p_Result_938_fu_10541_p3);

assign overflow_375_fu_10655_p2 = (xor_ln895_564_fu_10649_p2 & p_Result_940_fu_10641_p3);

assign overflow_fu_4056_p2 = (xor_ln895_485_fu_4051_p2 & or_ln895_fu_4046_p2);

assign p_Result_835_fu_5119_p3 = p_Val2_834_fu_5109_p2[32'd17];

assign p_Result_838_fu_5268_p3 = p_Val2_837_fu_5258_p2[32'd19];

assign p_Result_841_fu_5417_p3 = p_Val2_840_fu_5407_p2[32'd21];

assign p_Result_844_fu_5566_p3 = p_Val2_843_fu_5556_p2[32'd19];

assign p_Result_847_fu_5715_p3 = p_Val2_846_fu_5705_p2[32'd30];

assign p_Result_850_fu_5864_p3 = p_Val2_849_fu_5854_p2[32'd19];

assign p_Result_853_fu_6013_p3 = p_Val2_852_fu_6003_p2[32'd19];

assign p_Result_856_fu_6162_p3 = p_Val2_855_fu_6152_p2[32'd30];

assign p_Result_859_fu_6311_p3 = p_Val2_858_fu_6301_p2[32'd30];

assign p_Result_862_fu_8622_p3 = p_Val2_861_fu_8612_p2[32'd19];

assign p_Result_865_fu_8771_p3 = p_Val2_864_fu_8761_p2[32'd18];

assign p_Result_868_fu_8920_p3 = p_Val2_867_fu_8910_p2[32'd20];

assign p_Result_871_fu_9069_p3 = p_Val2_870_fu_9059_p2[32'd21];

assign p_Result_874_fu_9218_p3 = p_Val2_873_fu_9208_p2[32'd30];

assign p_Result_875_fu_3796_p3 = r_V_200_fu_3790_p2[32'd38];

assign p_Result_876_fu_3824_p3 = r_V_200_fu_3790_p2[32'd38];

assign p_Result_877_fu_3850_p3 = p_Val2_876_fu_3844_p2[32'd15];

assign p_Result_880_fu_9384_p3 = p_Val2_879_fu_9374_p2[32'd17];

assign p_Result_883_fu_9533_p3 = p_Val2_882_fu_9523_p2[32'd30];

assign p_Result_886_fu_9682_p3 = p_Val2_885_fu_9672_p2[32'd30];

assign p_Result_887_fu_6816_p3 = ret_V_fu_6810_p2[32'd32];

assign p_Result_888_fu_6830_p3 = p_Val2_887_fu_6824_p2[32'd31];

assign p_Result_889_fu_6914_p3 = ret_V_161_fu_6908_p2[32'd32];

assign p_Result_890_fu_6928_p3 = p_Val2_889_fu_6922_p2[32'd31];

assign p_Result_891_fu_7012_p3 = ret_V_162_fu_7006_p2[32'd32];

assign p_Result_892_fu_7026_p3 = p_Val2_891_fu_7020_p2[32'd31];

assign p_Result_893_fu_7110_p3 = ret_V_163_fu_7104_p2[32'd32];

assign p_Result_894_fu_7124_p3 = p_Val2_893_fu_7118_p2[32'd31];

assign p_Result_895_fu_7208_p3 = ret_V_164_fu_7202_p2[32'd32];

assign p_Result_896_fu_7222_p3 = p_Val2_895_fu_7216_p2[32'd31];

assign p_Result_897_fu_7306_p3 = ret_V_165_fu_7300_p2[32'd32];

assign p_Result_898_fu_7320_p3 = p_Val2_897_fu_7314_p2[32'd31];

assign p_Result_899_fu_7404_p3 = ret_V_166_fu_7398_p2[32'd32];

assign p_Result_900_fu_7418_p3 = p_Val2_899_fu_7412_p2[32'd31];

assign p_Result_901_fu_7502_p3 = ret_V_167_fu_7496_p2[32'd32];

assign p_Result_902_fu_7516_p3 = p_Val2_901_fu_7510_p2[32'd31];

assign p_Result_903_fu_7600_p3 = ret_V_168_fu_7594_p2[32'd32];

assign p_Result_904_fu_7614_p3 = p_Val2_903_fu_7608_p2[32'd31];

assign p_Result_905_fu_7702_p3 = ret_V_169_fu_7696_p2[32'd32];

assign p_Result_906_fu_7716_p3 = p_Val2_905_fu_7710_p2[32'd31];

assign p_Result_907_fu_7804_p3 = ret_V_170_fu_7798_p2[32'd32];

assign p_Result_908_fu_7818_p3 = p_Val2_907_fu_7812_p2[32'd31];

assign p_Result_909_fu_7906_p3 = ret_V_171_fu_7900_p2[32'd32];

assign p_Result_910_fu_7920_p3 = p_Val2_909_fu_7914_p2[32'd31];

assign p_Result_911_fu_8008_p3 = ret_V_172_fu_8002_p2[32'd32];

assign p_Result_912_fu_8022_p3 = p_Val2_911_fu_8016_p2[32'd31];

assign p_Result_913_fu_8110_p3 = ret_V_173_fu_8104_p2[32'd32];

assign p_Result_914_fu_8124_p3 = p_Val2_913_fu_8118_p2[32'd31];

assign p_Result_915_fu_8212_p3 = ret_V_174_fu_8206_p2[32'd32];

assign p_Result_916_fu_8226_p3 = p_Val2_915_fu_8220_p2[32'd31];

assign p_Result_917_fu_8314_p3 = ret_V_175_fu_8308_p2[32'd32];

assign p_Result_918_fu_8328_p3 = p_Val2_917_fu_8322_p2[32'd31];

assign p_Result_919_fu_8416_p3 = ret_V_176_fu_8410_p2[32'd32];

assign p_Result_920_fu_8430_p3 = p_Val2_919_fu_8424_p2[32'd31];

assign p_Result_921_fu_8518_p3 = ret_V_177_fu_8512_p2[32'd32];

assign p_Result_922_fu_8532_p3 = p_Val2_921_fu_8526_p2[32'd31];

assign p_Result_923_fu_9828_p3 = ret_V_178_fu_9822_p2[32'd32];

assign p_Result_924_fu_9841_p3 = p_Val2_923_fu_9836_p2[32'd31];

assign p_Result_925_fu_9928_p3 = ret_V_179_fu_9922_p2[32'd32];

assign p_Result_926_fu_9941_p3 = p_Val2_925_fu_9936_p2[32'd31];

assign p_Result_927_fu_10028_p3 = ret_V_180_fu_10022_p2[32'd32];

assign p_Result_928_fu_10041_p3 = p_Val2_927_fu_10036_p2[32'd31];

assign p_Result_929_fu_10128_p3 = ret_V_181_fu_10122_p2[32'd32];

assign p_Result_930_fu_10141_p3 = p_Val2_929_fu_10136_p2[32'd31];

assign p_Result_931_fu_10228_p3 = ret_V_182_fu_10222_p2[32'd32];

assign p_Result_932_fu_10241_p3 = p_Val2_931_fu_10236_p2[32'd31];

assign p_Result_933_fu_10328_p3 = ret_V_183_fu_10322_p2[32'd32];

assign p_Result_934_fu_10341_p3 = p_Val2_933_fu_10336_p2[32'd31];

assign p_Result_935_fu_10428_p3 = ret_V_184_fu_10422_p2[32'd32];

assign p_Result_936_fu_10441_p3 = p_Val2_935_fu_10436_p2[32'd31];

assign p_Result_937_fu_10528_p3 = ret_V_185_fu_10522_p2[32'd32];

assign p_Result_938_fu_10541_p3 = p_Val2_937_fu_10536_p2[32'd31];

assign p_Result_939_fu_10628_p3 = ret_V_186_fu_10622_p2[32'd32];

assign p_Result_940_fu_10641_p3 = p_Val2_939_fu_10636_p2[32'd31];

assign p_Val2_806_fu_2749_p4 = {{r_V_178_fu_254_p2[42:24]}};

assign p_Val2_807_fu_2783_p2 = ($signed(zext_ln377_fu_2779_p1) + $signed(sext_ln823_fu_2759_p1));

assign p_Val2_809_fu_2813_p4 = {{r_V_179_fu_262_p2[43:24]}};

assign p_Val2_810_fu_2847_p2 = ($signed(zext_ln377_161_fu_2843_p1) + $signed(sext_ln823_153_fu_2823_p1));

assign p_Val2_812_fu_2877_p4 = {{r_V_180_fu_251_p2[55:24]}};

assign p_Val2_813_fu_2907_p2 = (zext_ln377_162_fu_2903_p1 + p_Val2_812_fu_2877_p4);

assign p_Val2_815_fu_2937_p4 = {{r_V_181_fu_256_p2[43:24]}};

assign p_Val2_816_fu_2971_p2 = ($signed(zext_ln377_163_fu_2967_p1) + $signed(sext_ln823_154_fu_2947_p1));

assign p_Val2_818_fu_3001_p4 = {{r_V_182_fu_264_p2[46:24]}};

assign p_Val2_819_fu_3035_p2 = ($signed(zext_ln377_164_fu_3031_p1) + $signed(sext_ln823_155_fu_3011_p1));

assign p_Val2_821_fu_3065_p4 = {{r_V_183_fu_240_p2[42:24]}};

assign p_Val2_822_fu_3099_p2 = ($signed(zext_ln377_165_fu_3095_p1) + $signed(sext_ln823_156_fu_3075_p1));

assign p_Val2_824_fu_3129_p4 = {{r_V_184_fu_249_p2[42:24]}};

assign p_Val2_825_fu_3163_p2 = ($signed(zext_ln377_166_fu_3159_p1) + $signed(sext_ln823_157_fu_3139_p1));

assign p_Val2_827_fu_3193_p4 = {{r_V_185_fu_259_p2[53:24]}};

assign p_Val2_828_fu_3227_p2 = ($signed(zext_ln377_167_fu_3223_p1) + $signed(sext_ln823_158_fu_3203_p1));

assign p_Val2_830_fu_3257_p4 = {{r_V_186_fu_246_p2[53:24]}};

assign p_Val2_831_fu_3291_p2 = ($signed(zext_ln377_168_fu_3287_p1) + $signed(sext_ln823_159_fu_3267_p1));

assign p_Val2_834_fu_5109_p2 = ($signed(zext_ln377_169_fu_5106_p1) + $signed(sext_ln823_160_fu_5103_p1));

assign p_Val2_837_fu_5258_p2 = ($signed(zext_ln377_170_fu_5255_p1) + $signed(sext_ln823_161_fu_5252_p1));

assign p_Val2_840_fu_5407_p2 = ($signed(zext_ln377_171_fu_5404_p1) + $signed(sext_ln823_162_fu_5401_p1));

assign p_Val2_843_fu_5556_p2 = ($signed(zext_ln377_172_fu_5553_p1) + $signed(sext_ln823_163_fu_5550_p1));

assign p_Val2_846_fu_5705_p2 = ($signed(zext_ln377_173_fu_5702_p1) + $signed(sext_ln823_164_fu_5699_p1));

assign p_Val2_849_fu_5854_p2 = ($signed(zext_ln377_174_fu_5851_p1) + $signed(sext_ln823_165_fu_5848_p1));

assign p_Val2_852_fu_6003_p2 = ($signed(zext_ln377_175_fu_6000_p1) + $signed(sext_ln823_166_fu_5997_p1));

assign p_Val2_855_fu_6152_p2 = ($signed(zext_ln377_176_fu_6149_p1) + $signed(sext_ln823_167_fu_6146_p1));

assign p_Val2_858_fu_6301_p2 = ($signed(zext_ln377_177_fu_6298_p1) + $signed(sext_ln823_168_fu_6295_p1));

assign p_Val2_861_fu_8612_p2 = ($signed(zext_ln377_178_fu_8609_p1) + $signed(sext_ln823_169_fu_8606_p1));

assign p_Val2_864_fu_8761_p2 = ($signed(zext_ln377_179_fu_8758_p1) + $signed(sext_ln823_170_fu_8755_p1));

assign p_Val2_867_fu_8910_p2 = ($signed(zext_ln377_180_fu_8907_p1) + $signed(sext_ln823_171_fu_8904_p1));

assign p_Val2_870_fu_9059_p2 = ($signed(zext_ln377_181_fu_9056_p1) + $signed(sext_ln823_172_fu_9053_p1));

assign p_Val2_873_fu_9208_p2 = ($signed(zext_ln377_182_fu_9205_p1) + $signed(sext_ln823_173_fu_9202_p1));

assign p_Val2_875_fu_3804_p4 = {{r_V_200_fu_3790_p2[38:24]}};

assign p_Val2_876_fu_3844_p2 = ($signed(zext_ln377_183_fu_3840_p1) + $signed(sext_ln823_174_fu_3814_p1));

assign p_Val2_879_fu_9374_p2 = ($signed(zext_ln377_184_fu_9371_p1) + $signed(sext_ln823_175_fu_9368_p1));

assign p_Val2_882_fu_9523_p2 = ($signed(zext_ln377_185_fu_9520_p1) + $signed(sext_ln823_176_fu_9517_p1));

assign p_Val2_885_fu_9672_p2 = ($signed(zext_ln377_186_fu_9669_p1) + $signed(sext_ln823_177_fu_9666_p1));

assign p_Val2_887_fu_6824_p2 = ($signed(rhs_fu_4099_p3) + $signed(32'd4294960969));

assign p_Val2_889_fu_6922_p2 = ($signed(rhs_161_fu_4224_p3) + $signed(32'd4294801704));

assign p_Val2_891_fu_7020_p2 = ($signed(rhs_162_fu_4346_p3) + $signed(32'd4294057118));

assign p_Val2_893_fu_7118_p2 = ($signed(rhs_163_fu_4470_p3) + $signed(32'd4294941217));

assign p_Val2_895_fu_7216_p2 = ($signed(rhs_164_fu_4595_p3) + $signed(32'd5765636));

assign p_Val2_897_fu_7314_p2 = ($signed(rhs_165_fu_4720_p3) + $signed(32'd4294963905));

assign p_Val2_899_fu_7412_p2 = ($signed(rhs_166_fu_4845_p3) + $signed(32'd4294962962));

assign p_Val2_901_fu_7510_p2 = ($signed(rhs_167_fu_4970_p3) + $signed(32'd4294697172));

assign p_Val2_903_fu_7608_p2 = ($signed(rhs_168_fu_5095_p3) + $signed(32'd4293009208));

assign p_Val2_905_fu_7710_p2 = ($signed(rhs_169_fu_5244_p3) + $signed(lhs_fu_6896_p3));

assign p_Val2_907_fu_7812_p2 = ($signed(rhs_170_fu_5393_p3) + $signed(lhs_143_fu_6994_p3));

assign p_Val2_909_fu_7914_p2 = ($signed(rhs_171_fu_5542_p3) + $signed(lhs_144_fu_7092_p3));

assign p_Val2_911_fu_8016_p2 = ($signed(rhs_172_fu_5691_p3) + $signed(lhs_145_fu_7190_p3));

assign p_Val2_913_fu_8118_p2 = ($signed(rhs_173_fu_5840_p3) + $signed(lhs_146_fu_7288_p3));

assign p_Val2_915_fu_8220_p2 = ($signed(rhs_174_fu_5989_p3) + $signed(lhs_147_fu_7386_p3));

assign p_Val2_917_fu_8322_p2 = ($signed(rhs_175_fu_6138_p3) + $signed(lhs_148_fu_7484_p3));

assign p_Val2_919_fu_8424_p2 = ($signed(rhs_176_fu_6287_p3) + $signed(lhs_149_fu_7582_p3));

assign p_Val2_921_fu_8526_p2 = ($signed(rhs_177_fu_6436_p3) + $signed(lhs_150_fu_7680_p3));

assign p_Val2_923_fu_9836_p2 = ($signed(rhs_178_fu_8747_p3) + $signed(lhs_151_reg_11566));

assign p_Val2_925_fu_9936_p2 = ($signed(rhs_179_fu_8896_p3) + $signed(lhs_152_reg_11572));

assign p_Val2_927_fu_10036_p2 = ($signed(rhs_180_fu_9045_p3) + $signed(lhs_153_reg_11578));

assign p_Val2_929_fu_10136_p2 = ($signed(rhs_181_fu_9194_p3) + $signed(lhs_154_reg_11584));

assign p_Val2_931_fu_10236_p2 = ($signed(rhs_182_fu_9343_p3) + $signed(lhs_155_reg_11590));

assign p_Val2_933_fu_10336_p2 = ($signed(rhs_183_fu_9361_p3) + $signed(lhs_156_reg_11596));

assign p_Val2_935_fu_10436_p2 = ($signed(rhs_184_fu_9509_p3) + $signed(lhs_157_reg_11602));

assign p_Val2_937_fu_10536_p2 = ($signed(rhs_185_fu_9658_p3) + $signed(lhs_158_reg_11608));

assign p_Val2_939_fu_10636_p2 = ($signed(rhs_186_fu_9807_p3) + $signed(lhs_159_reg_11614));

assign r_V_178_fu_254_p0 = sext_ln70_93_fu_2734_p1;

assign r_V_178_fu_254_p1 = 43'd8796093021447;

assign r_V_179_fu_262_p0 = sext_ln70_92_fu_2728_p1;

assign r_V_179_fu_262_p1 = 44'd17592186043026;

assign r_V_180_fu_251_p1 = 57'd25766628;

assign r_V_181_fu_256_p0 = sext_ln70_92_fu_2728_p1;

assign r_V_181_fu_256_p1 = 44'd17592186043035;

assign r_V_182_fu_264_p1 = 47'd12067;

assign r_V_183_fu_240_p0 = sext_ln70_93_fu_2734_p1;

assign r_V_183_fu_240_p1 = 43'd558;

assign r_V_184_fu_249_p0 = sext_ln70_93_fu_2734_p1;

assign r_V_184_fu_249_p1 = 43'd901;

assign r_V_185_fu_259_p0 = sext_ln70_fu_2712_p1;

assign r_V_185_fu_259_p1 = 54'd2291250;

assign r_V_186_fu_246_p0 = sext_ln70_fu_2712_p1;

assign r_V_186_fu_246_p1 = 54'd2264876;

assign r_V_187_fu_266_p1 = 41'd2199023255395;

assign r_V_188_fu_261_p0 = sext_ln70_96_fu_3335_p1;

assign r_V_188_fu_261_p1 = 43'd805;

assign r_V_189_fu_242_p1 = 45'd35184372084910;

assign r_V_190_fu_260_p0 = sext_ln70_96_fu_3335_p1;

assign r_V_190_fu_260_p1 = 43'd525;

assign r_V_191_fu_263_p0 = sext_ln70_94_fu_3323_p1;

assign r_V_191_fu_263_p1 = 54'd3046284;

assign r_V_192_fu_250_p0 = sext_ln70_96_fu_3335_p1;

assign r_V_192_fu_250_p1 = 43'd860;

assign r_V_193_fu_244_p0 = sext_ln70_96_fu_3335_p1;

assign r_V_193_fu_244_p1 = 43'd8796093021252;

assign r_V_194_fu_243_p0 = sext_ln70_94_fu_3323_p1;

assign r_V_194_fu_243_p1 = 54'd18014398506808642;

assign r_V_195_fu_248_p0 = sext_ln70_94_fu_3323_p1;

assign r_V_195_fu_248_p1 = 54'd18014398506836554;

assign r_V_196_fu_258_p1 = 42'd4398046510642;

assign r_V_197_fu_245_p1 = 44'd1347;

assign r_V_198_fu_265_p1 = 45'd35184372086576;

assign r_V_199_fu_255_p0 = sext_ln70_100_fu_6448_p1;

assign r_V_199_fu_255_p1 = 54'd18014398506422962;

assign r_V_200_fu_3790_p2 = ($signed(sext_ln1273_fu_3768_p1) + $signed(sext_ln70_99_fu_3746_p1));

assign r_V_201_fu_257_p1 = 41'd2199023255347;

assign r_V_202_fu_252_p0 = sext_ln70_100_fu_6448_p1;

assign r_V_202_fu_252_p1 = 54'd2644459;

assign r_V_203_fu_253_p0 = sext_ln70_100_fu_6448_p1;

assign r_V_203_fu_253_p1 = 54'd2578651;

assign r_V_fu_247_p1 = 43'd8796093021602;

assign ret_V_161_fu_6908_p2 = ($signed(sext_ln813_305_fu_6904_p1) + $signed(33'd8589769000));

assign ret_V_162_fu_7006_p2 = ($signed(sext_ln813_306_fu_7002_p1) + $signed(33'd8589024414));

assign ret_V_163_fu_7104_p2 = ($signed(sext_ln813_307_fu_7100_p1) + $signed(33'd8589908513));

assign ret_V_164_fu_7202_p2 = ($signed(sext_ln813_308_fu_7198_p1) + $signed(33'd5765636));

assign ret_V_165_fu_7300_p2 = ($signed(sext_ln813_309_fu_7296_p1) + $signed(33'd8589931201));

assign ret_V_166_fu_7398_p2 = ($signed(sext_ln813_310_fu_7394_p1) + $signed(33'd8589930258));

assign ret_V_167_fu_7496_p2 = ($signed(sext_ln813_311_fu_7492_p1) + $signed(33'd8589664468));

assign ret_V_168_fu_7594_p2 = ($signed(sext_ln813_312_fu_7590_p1) + $signed(33'd8587976504));

assign ret_V_169_fu_7696_p2 = ($signed(sext_ln813_314_fu_7692_p1) + $signed(sext_ln813_313_fu_7688_p1));

assign ret_V_170_fu_7798_p2 = ($signed(sext_ln813_316_fu_7794_p1) + $signed(sext_ln813_315_fu_7790_p1));

assign ret_V_171_fu_7900_p2 = ($signed(sext_ln813_318_fu_7896_p1) + $signed(sext_ln813_317_fu_7892_p1));

assign ret_V_172_fu_8002_p2 = ($signed(sext_ln813_320_fu_7998_p1) + $signed(sext_ln813_319_fu_7994_p1));

assign ret_V_173_fu_8104_p2 = ($signed(sext_ln813_322_fu_8100_p1) + $signed(sext_ln813_321_fu_8096_p1));

assign ret_V_174_fu_8206_p2 = ($signed(sext_ln813_324_fu_8202_p1) + $signed(sext_ln813_323_fu_8198_p1));

assign ret_V_175_fu_8308_p2 = ($signed(sext_ln813_326_fu_8304_p1) + $signed(sext_ln813_325_fu_8300_p1));

assign ret_V_176_fu_8410_p2 = ($signed(sext_ln813_328_fu_8406_p1) + $signed(sext_ln813_327_fu_8402_p1));

assign ret_V_177_fu_8512_p2 = ($signed(sext_ln813_330_fu_8508_p1) + $signed(sext_ln813_329_fu_8504_p1));

assign ret_V_178_fu_9822_p2 = ($signed(sext_ln813_332_fu_9818_p1) + $signed(sext_ln813_331_fu_9815_p1));

assign ret_V_179_fu_9922_p2 = ($signed(sext_ln813_334_fu_9918_p1) + $signed(sext_ln813_333_fu_9915_p1));

assign ret_V_180_fu_10022_p2 = ($signed(sext_ln813_336_fu_10018_p1) + $signed(sext_ln813_335_fu_10015_p1));

assign ret_V_181_fu_10122_p2 = ($signed(sext_ln813_338_fu_10118_p1) + $signed(sext_ln813_337_fu_10115_p1));

assign ret_V_182_fu_10222_p2 = ($signed(sext_ln813_340_fu_10218_p1) + $signed(sext_ln813_339_fu_10215_p1));

assign ret_V_183_fu_10322_p2 = ($signed(sext_ln813_342_fu_10318_p1) + $signed(sext_ln813_341_fu_10315_p1));

assign ret_V_184_fu_10422_p2 = ($signed(sext_ln813_344_fu_10418_p1) + $signed(sext_ln813_343_fu_10415_p1));

assign ret_V_185_fu_10522_p2 = ($signed(sext_ln813_346_fu_10518_p1) + $signed(sext_ln813_345_fu_10515_p1));

assign ret_V_186_fu_10622_p2 = ($signed(sext_ln813_348_fu_10618_p1) + $signed(sext_ln813_347_fu_10615_p1));

assign ret_V_fu_6810_p2 = ($signed(sext_ln813_fu_6806_p1) + $signed(33'd8589928265));

assign rhs_161_fu_4224_p3 = ((or_ln346_161_fu_4218_p2[0:0] == 1'b1) ? select_ln346_244_fu_4210_p3 : sext_ln856_153_fu_4107_p1);

assign rhs_162_fu_4346_p3 = ((or_ln346_162_fu_4340_p2[0:0] == 1'b1) ? select_ln346_245_fu_4332_p3 : p_Val2_813_reg_10843);

assign rhs_163_fu_4470_p3 = ((or_ln346_163_fu_4464_p2[0:0] == 1'b1) ? select_ln346_246_fu_4456_p3 : sext_ln856_154_fu_4353_p1);

assign rhs_164_fu_4595_p3 = ((or_ln346_164_fu_4589_p2[0:0] == 1'b1) ? select_ln346_247_fu_4581_p3 : sext_ln856_155_fu_4478_p1);

assign rhs_165_fu_4720_p3 = ((or_ln346_165_fu_4714_p2[0:0] == 1'b1) ? select_ln346_248_fu_4706_p3 : sext_ln856_156_fu_4603_p1);

assign rhs_166_fu_4845_p3 = ((or_ln346_166_fu_4839_p2[0:0] == 1'b1) ? select_ln346_249_fu_4831_p3 : sext_ln856_157_fu_4728_p1);

assign rhs_167_fu_4970_p3 = ((or_ln346_167_fu_4964_p2[0:0] == 1'b1) ? select_ln346_250_fu_4956_p3 : sext_ln856_158_fu_4853_p1);

assign rhs_168_fu_5095_p3 = ((or_ln346_168_fu_5089_p2[0:0] == 1'b1) ? select_ln346_251_fu_5081_p3 : sext_ln856_159_fu_4978_p1);

assign rhs_169_fu_5244_p3 = ((or_ln346_169_fu_5238_p2[0:0] == 1'b1) ? select_ln346_252_fu_5230_p3 : sext_ln856_160_fu_5115_p1);

assign rhs_170_fu_5393_p3 = ((or_ln346_170_fu_5387_p2[0:0] == 1'b1) ? select_ln346_253_fu_5379_p3 : sext_ln856_161_fu_5264_p1);

assign rhs_171_fu_5542_p3 = ((or_ln346_171_fu_5536_p2[0:0] == 1'b1) ? select_ln346_254_fu_5528_p3 : sext_ln856_162_fu_5413_p1);

assign rhs_172_fu_5691_p3 = ((or_ln346_172_fu_5685_p2[0:0] == 1'b1) ? select_ln346_255_fu_5677_p3 : sext_ln856_163_fu_5562_p1);

assign rhs_173_fu_5840_p3 = ((or_ln346_173_fu_5834_p2[0:0] == 1'b1) ? select_ln346_256_fu_5826_p3 : sext_ln856_164_fu_5711_p1);

assign rhs_174_fu_5989_p3 = ((or_ln346_174_fu_5983_p2[0:0] == 1'b1) ? select_ln346_257_fu_5975_p3 : sext_ln856_165_fu_5860_p1);

assign rhs_175_fu_6138_p3 = ((or_ln346_175_fu_6132_p2[0:0] == 1'b1) ? select_ln346_258_fu_6124_p3 : sext_ln856_166_fu_6009_p1);

assign rhs_176_fu_6287_p3 = ((or_ln346_176_fu_6281_p2[0:0] == 1'b1) ? select_ln346_259_fu_6273_p3 : sext_ln856_167_fu_6158_p1);

assign rhs_177_fu_6436_p3 = ((or_ln346_177_fu_6430_p2[0:0] == 1'b1) ? select_ln346_260_fu_6422_p3 : sext_ln856_168_fu_6307_p1);

assign rhs_178_fu_8747_p3 = ((or_ln346_178_fu_8741_p2[0:0] == 1'b1) ? select_ln346_261_fu_8733_p3 : sext_ln856_169_fu_8618_p1);

assign rhs_179_fu_8896_p3 = ((or_ln346_179_fu_8890_p2[0:0] == 1'b1) ? select_ln346_262_fu_8882_p3 : sext_ln856_170_fu_8767_p1);

assign rhs_180_fu_9045_p3 = ((or_ln346_180_fu_9039_p2[0:0] == 1'b1) ? select_ln346_263_fu_9031_p3 : sext_ln856_171_fu_8916_p1);

assign rhs_181_fu_9194_p3 = ((or_ln346_181_fu_9188_p2[0:0] == 1'b1) ? select_ln346_264_fu_9180_p3 : sext_ln856_172_fu_9065_p1);

assign rhs_182_fu_9343_p3 = ((or_ln346_182_fu_9337_p2[0:0] == 1'b1) ? select_ln346_265_fu_9329_p3 : sext_ln856_173_fu_9214_p1);

assign rhs_183_fu_9361_p3 = ((or_ln346_183_reg_11329_pp0_iter1_reg[0:0] == 1'b1) ? select_ln346_266_fu_9354_p3 : sext_ln856_174_fu_9351_p1);

assign rhs_184_fu_9509_p3 = ((or_ln346_184_fu_9503_p2[0:0] == 1'b1) ? select_ln346_267_fu_9495_p3 : sext_ln856_175_fu_9380_p1);

assign rhs_185_fu_9658_p3 = ((or_ln346_185_fu_9652_p2[0:0] == 1'b1) ? select_ln346_268_fu_9644_p3 : sext_ln856_176_fu_9529_p1);

assign rhs_186_fu_9807_p3 = ((or_ln346_186_fu_9801_p2[0:0] == 1'b1) ? select_ln346_269_fu_9793_p3 : sext_ln856_177_fu_9678_p1);

assign rhs_fu_4099_p3 = ((or_ln346_fu_4093_p2[0:0] == 1'b1) ? select_ln346_243_fu_4085_p3 : sext_ln856_fu_3982_p1);

assign select_ln302_324_fu_6978_p3 = ((xor_ln302_324_fu_6960_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_889_fu_6922_p2);

assign select_ln302_326_fu_7076_p3 = ((xor_ln302_326_fu_7058_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_891_fu_7020_p2);

assign select_ln302_328_fu_7174_p3 = ((xor_ln302_328_fu_7156_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_893_fu_7118_p2);

assign select_ln302_330_fu_7272_p3 = ((xor_ln302_330_fu_7254_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_895_fu_7216_p2);

assign select_ln302_332_fu_7370_p3 = ((xor_ln302_332_fu_7352_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_897_fu_7314_p2);

assign select_ln302_334_fu_7468_p3 = ((xor_ln302_334_fu_7450_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_899_fu_7412_p2);

assign select_ln302_336_fu_7566_p3 = ((xor_ln302_336_fu_7548_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_901_fu_7510_p2);

assign select_ln302_338_fu_7664_p3 = ((xor_ln302_338_fu_7646_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_903_fu_7608_p2);

assign select_ln302_340_fu_7766_p3 = ((xor_ln302_340_fu_7748_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_905_fu_7710_p2);

assign select_ln302_342_fu_7868_p3 = ((xor_ln302_342_fu_7850_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_907_fu_7812_p2);

assign select_ln302_344_fu_7970_p3 = ((xor_ln302_344_fu_7952_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_909_fu_7914_p2);

assign select_ln302_346_fu_8072_p3 = ((xor_ln302_346_fu_8054_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_911_fu_8016_p2);

assign select_ln302_348_fu_8174_p3 = ((xor_ln302_348_fu_8156_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_913_fu_8118_p2);

assign select_ln302_350_fu_8276_p3 = ((xor_ln302_350_fu_8258_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_915_fu_8220_p2);

assign select_ln302_352_fu_8378_p3 = ((xor_ln302_352_fu_8360_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_917_fu_8322_p2);

assign select_ln302_354_fu_8480_p3 = ((xor_ln302_354_fu_8462_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_919_fu_8424_p2);

assign select_ln302_356_fu_8582_p3 = ((xor_ln302_356_fu_8564_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_921_fu_8526_p2);

assign select_ln302_358_fu_9891_p3 = ((xor_ln302_358_fu_9873_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_923_fu_9836_p2);

assign select_ln302_359_fu_9907_p3 = ((or_ln302_178_fu_9885_p2[0:0] == 1'b1) ? select_ln302_358_fu_9891_p3 : select_ln350_178_fu_9899_p3);

assign select_ln302_360_fu_9991_p3 = ((xor_ln302_360_fu_9973_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_925_fu_9936_p2);

assign select_ln302_361_fu_10007_p3 = ((or_ln302_179_fu_9985_p2[0:0] == 1'b1) ? select_ln302_360_fu_9991_p3 : select_ln350_179_fu_9999_p3);

assign select_ln302_362_fu_10091_p3 = ((xor_ln302_362_fu_10073_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_927_fu_10036_p2);

assign select_ln302_363_fu_10107_p3 = ((or_ln302_180_fu_10085_p2[0:0] == 1'b1) ? select_ln302_362_fu_10091_p3 : select_ln350_180_fu_10099_p3);

assign select_ln302_364_fu_10191_p3 = ((xor_ln302_364_fu_10173_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_929_fu_10136_p2);

assign select_ln302_365_fu_10207_p3 = ((or_ln302_181_fu_10185_p2[0:0] == 1'b1) ? select_ln302_364_fu_10191_p3 : select_ln350_181_fu_10199_p3);

assign select_ln302_366_fu_10291_p3 = ((xor_ln302_366_fu_10273_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_931_fu_10236_p2);

assign select_ln302_367_fu_10307_p3 = ((or_ln302_182_fu_10285_p2[0:0] == 1'b1) ? select_ln302_366_fu_10291_p3 : select_ln350_182_fu_10299_p3);

assign select_ln302_368_fu_10391_p3 = ((xor_ln302_368_fu_10373_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_933_fu_10336_p2);

assign select_ln302_369_fu_10407_p3 = ((or_ln302_183_fu_10385_p2[0:0] == 1'b1) ? select_ln302_368_fu_10391_p3 : select_ln350_183_fu_10399_p3);

assign select_ln302_370_fu_10491_p3 = ((xor_ln302_370_fu_10473_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_935_fu_10436_p2);

assign select_ln302_371_fu_10507_p3 = ((or_ln302_184_fu_10485_p2[0:0] == 1'b1) ? select_ln302_370_fu_10491_p3 : select_ln350_184_fu_10499_p3);

assign select_ln302_372_fu_10591_p3 = ((xor_ln302_372_fu_10573_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_937_fu_10536_p2);

assign select_ln302_373_fu_10607_p3 = ((or_ln302_185_fu_10585_p2[0:0] == 1'b1) ? select_ln302_372_fu_10591_p3 : select_ln350_185_fu_10599_p3);

assign select_ln302_374_fu_10691_p3 = ((xor_ln302_374_fu_10673_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_939_fu_10636_p2);

assign select_ln302_375_fu_10707_p3 = ((or_ln302_186_fu_10685_p2[0:0] == 1'b1) ? select_ln302_374_fu_10691_p3 : select_ln350_186_fu_10699_p3);

assign select_ln302_fu_6880_p3 = ((xor_ln302_fu_6862_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_887_fu_6824_p2);

assign select_ln346_243_fu_4085_p3 = ((overflow_fu_4056_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_244_fu_4210_p3 = ((overflow_323_fu_4181_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_245_fu_4332_p3 = ((overflow_324_fu_4303_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_246_fu_4456_p3 = ((overflow_325_fu_4427_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_247_fu_4581_p3 = ((overflow_326_fu_4552_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_248_fu_4706_p3 = ((overflow_327_fu_4677_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_249_fu_4831_p3 = ((overflow_328_fu_4802_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_250_fu_4956_p3 = ((overflow_329_fu_4927_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_251_fu_5081_p3 = ((overflow_330_fu_5052_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_252_fu_5230_p3 = ((overflow_331_fu_5201_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_253_fu_5379_p3 = ((overflow_332_fu_5350_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_254_fu_5528_p3 = ((overflow_333_fu_5499_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_255_fu_5677_p3 = ((overflow_334_fu_5648_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_256_fu_5826_p3 = ((overflow_335_fu_5797_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_257_fu_5975_p3 = ((overflow_336_fu_5946_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_258_fu_6124_p3 = ((overflow_337_fu_6095_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_259_fu_6273_p3 = ((overflow_338_fu_6244_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_260_fu_6422_p3 = ((overflow_339_fu_6393_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_261_fu_8733_p3 = ((overflow_340_fu_8704_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_262_fu_8882_p3 = ((overflow_341_fu_8853_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_263_fu_9031_p3 = ((overflow_342_fu_9002_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_264_fu_9180_p3 = ((overflow_343_fu_9151_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_265_fu_9329_p3 = ((overflow_344_fu_9300_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_266_fu_9354_p3 = ((overflow_345_reg_11324_pp0_iter1_reg[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_267_fu_9495_p3 = ((overflow_346_fu_9466_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_268_fu_9644_p3 = ((overflow_347_fu_9615_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_269_fu_9793_p3 = ((overflow_348_fu_9764_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln350_161_fu_6986_p3 = ((underflow_350_fu_6954_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_889_fu_6922_p2);

assign select_ln350_162_fu_7084_p3 = ((underflow_351_fu_7052_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_891_fu_7020_p2);

assign select_ln350_163_fu_7182_p3 = ((underflow_352_fu_7150_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_893_fu_7118_p2);

assign select_ln350_164_fu_7280_p3 = ((underflow_353_fu_7248_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_895_fu_7216_p2);

assign select_ln350_165_fu_7378_p3 = ((underflow_354_fu_7346_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_897_fu_7314_p2);

assign select_ln350_166_fu_7476_p3 = ((underflow_355_fu_7444_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_899_fu_7412_p2);

assign select_ln350_167_fu_7574_p3 = ((underflow_356_fu_7542_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_901_fu_7510_p2);

assign select_ln350_168_fu_7672_p3 = ((underflow_357_fu_7640_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_903_fu_7608_p2);

assign select_ln350_169_fu_7774_p3 = ((underflow_358_fu_7742_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_905_fu_7710_p2);

assign select_ln350_170_fu_7876_p3 = ((underflow_359_fu_7844_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_907_fu_7812_p2);

assign select_ln350_171_fu_7978_p3 = ((underflow_360_fu_7946_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_909_fu_7914_p2);

assign select_ln350_172_fu_8080_p3 = ((underflow_361_fu_8048_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_911_fu_8016_p2);

assign select_ln350_173_fu_8182_p3 = ((underflow_362_fu_8150_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_913_fu_8118_p2);

assign select_ln350_174_fu_8284_p3 = ((underflow_363_fu_8252_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_915_fu_8220_p2);

assign select_ln350_175_fu_8386_p3 = ((underflow_364_fu_8354_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_917_fu_8322_p2);

assign select_ln350_176_fu_8488_p3 = ((underflow_365_fu_8456_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_919_fu_8424_p2);

assign select_ln350_177_fu_8590_p3 = ((underflow_366_fu_8558_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_921_fu_8526_p2);

assign select_ln350_178_fu_9899_p3 = ((underflow_367_fu_9867_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_923_fu_9836_p2);

assign select_ln350_179_fu_9999_p3 = ((underflow_368_fu_9967_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_925_fu_9936_p2);

assign select_ln350_180_fu_10099_p3 = ((underflow_369_fu_10067_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_927_fu_10036_p2);

assign select_ln350_181_fu_10199_p3 = ((underflow_370_fu_10167_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_929_fu_10136_p2);

assign select_ln350_182_fu_10299_p3 = ((underflow_371_fu_10267_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_931_fu_10236_p2);

assign select_ln350_183_fu_10399_p3 = ((underflow_372_fu_10367_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_933_fu_10336_p2);

assign select_ln350_184_fu_10499_p3 = ((underflow_373_fu_10467_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_935_fu_10436_p2);

assign select_ln350_185_fu_10599_p3 = ((underflow_374_fu_10567_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_937_fu_10536_p2);

assign select_ln350_186_fu_10699_p3 = ((underflow_375_fu_10667_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_939_fu_10636_p2);

assign select_ln350_fu_6888_p3 = ((underflow_349_fu_6856_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_887_fu_6824_p2);

assign sext_ln1273_fu_3768_p1 = $signed(shl_ln_fu_3760_p3);

assign sext_ln70_100_fu_6448_p1 = a_V_2_reg_11309;

assign sext_ln70_92_fu_2728_p1 = a_V_fu_2708_p1;

assign sext_ln70_93_fu_2734_p1 = a_V_fu_2708_p1;

assign sext_ln70_94_fu_3323_p1 = a_V_1_fu_3313_p4;

assign sext_ln70_96_fu_3335_p1 = a_V_1_fu_3313_p4;

assign sext_ln70_99_fu_3746_p1 = a_V_2_fu_3726_p4;

assign sext_ln70_fu_2712_p1 = a_V_fu_2708_p1;

assign sext_ln813_305_fu_6904_p1 = rhs_161_fu_4224_p3;

assign sext_ln813_306_fu_7002_p1 = rhs_162_fu_4346_p3;

assign sext_ln813_307_fu_7100_p1 = rhs_163_fu_4470_p3;

assign sext_ln813_308_fu_7198_p1 = rhs_164_fu_4595_p3;

assign sext_ln813_309_fu_7296_p1 = rhs_165_fu_4720_p3;

assign sext_ln813_310_fu_7394_p1 = rhs_166_fu_4845_p3;

assign sext_ln813_311_fu_7492_p1 = rhs_167_fu_4970_p3;

assign sext_ln813_312_fu_7590_p1 = rhs_168_fu_5095_p3;

assign sext_ln813_313_fu_7688_p1 = lhs_fu_6896_p3;

assign sext_ln813_314_fu_7692_p1 = rhs_169_fu_5244_p3;

assign sext_ln813_315_fu_7790_p1 = lhs_143_fu_6994_p3;

assign sext_ln813_316_fu_7794_p1 = rhs_170_fu_5393_p3;

assign sext_ln813_317_fu_7892_p1 = lhs_144_fu_7092_p3;

assign sext_ln813_318_fu_7896_p1 = rhs_171_fu_5542_p3;

assign sext_ln813_319_fu_7994_p1 = lhs_145_fu_7190_p3;

assign sext_ln813_320_fu_7998_p1 = rhs_172_fu_5691_p3;

assign sext_ln813_321_fu_8096_p1 = lhs_146_fu_7288_p3;

assign sext_ln813_322_fu_8100_p1 = rhs_173_fu_5840_p3;

assign sext_ln813_323_fu_8198_p1 = lhs_147_fu_7386_p3;

assign sext_ln813_324_fu_8202_p1 = rhs_174_fu_5989_p3;

assign sext_ln813_325_fu_8300_p1 = lhs_148_fu_7484_p3;

assign sext_ln813_326_fu_8304_p1 = rhs_175_fu_6138_p3;

assign sext_ln813_327_fu_8402_p1 = lhs_149_fu_7582_p3;

assign sext_ln813_328_fu_8406_p1 = rhs_176_fu_6287_p3;

assign sext_ln813_329_fu_8504_p1 = lhs_150_fu_7680_p3;

assign sext_ln813_330_fu_8508_p1 = rhs_177_fu_6436_p3;

assign sext_ln813_331_fu_9815_p1 = lhs_151_reg_11566;

assign sext_ln813_332_fu_9818_p1 = rhs_178_fu_8747_p3;

assign sext_ln813_333_fu_9915_p1 = lhs_152_reg_11572;

assign sext_ln813_334_fu_9918_p1 = rhs_179_fu_8896_p3;

assign sext_ln813_335_fu_10015_p1 = lhs_153_reg_11578;

assign sext_ln813_336_fu_10018_p1 = rhs_180_fu_9045_p3;

assign sext_ln813_337_fu_10115_p1 = lhs_154_reg_11584;

assign sext_ln813_338_fu_10118_p1 = rhs_181_fu_9194_p3;

assign sext_ln813_339_fu_10215_p1 = lhs_155_reg_11590;

assign sext_ln813_340_fu_10218_p1 = rhs_182_fu_9343_p3;

assign sext_ln813_341_fu_10315_p1 = lhs_156_reg_11596;

assign sext_ln813_342_fu_10318_p1 = rhs_183_fu_9361_p3;

assign sext_ln813_343_fu_10415_p1 = lhs_157_reg_11602;

assign sext_ln813_344_fu_10418_p1 = rhs_184_fu_9509_p3;

assign sext_ln813_345_fu_10515_p1 = lhs_158_reg_11608;

assign sext_ln813_346_fu_10518_p1 = rhs_185_fu_9658_p3;

assign sext_ln813_347_fu_10615_p1 = lhs_159_reg_11614;

assign sext_ln813_348_fu_10618_p1 = rhs_186_fu_9807_p3;

assign sext_ln813_fu_6806_p1 = rhs_fu_4099_p3;

assign sext_ln823_153_fu_2823_p1 = $signed(p_Val2_809_fu_2813_p4);

assign sext_ln823_154_fu_2947_p1 = $signed(p_Val2_815_fu_2937_p4);

assign sext_ln823_155_fu_3011_p1 = $signed(p_Val2_818_fu_3001_p4);

assign sext_ln823_156_fu_3075_p1 = $signed(p_Val2_821_fu_3065_p4);

assign sext_ln823_157_fu_3139_p1 = $signed(p_Val2_824_fu_3129_p4);

assign sext_ln823_158_fu_3203_p1 = $signed(p_Val2_827_fu_3193_p4);

assign sext_ln823_159_fu_3267_p1 = $signed(p_Val2_830_fu_3257_p4);

assign sext_ln823_160_fu_5103_p1 = $signed(p_Val2_833_reg_11054);

assign sext_ln823_161_fu_5252_p1 = $signed(p_Val2_836_reg_11083);

assign sext_ln823_162_fu_5401_p1 = $signed(p_Val2_839_reg_11112);

assign sext_ln823_163_fu_5550_p1 = $signed(p_Val2_842_reg_11141);

assign sext_ln823_164_fu_5699_p1 = $signed(p_Val2_845_reg_11170);

assign sext_ln823_165_fu_5848_p1 = $signed(p_Val2_848_reg_11199);

assign sext_ln823_166_fu_5997_p1 = $signed(p_Val2_851_reg_11228);

assign sext_ln823_167_fu_6146_p1 = $signed(p_Val2_854_reg_11257);

assign sext_ln823_168_fu_6295_p1 = $signed(p_Val2_857_reg_11286);

assign sext_ln823_169_fu_8606_p1 = $signed(p_Val2_860_reg_11340);

assign sext_ln823_170_fu_8755_p1 = $signed(p_Val2_863_reg_11369);

assign sext_ln823_171_fu_8904_p1 = $signed(p_Val2_866_reg_11398);

assign sext_ln823_172_fu_9053_p1 = $signed(p_Val2_869_reg_11427);

assign sext_ln823_173_fu_9202_p1 = $signed(p_Val2_872_reg_11456);

assign sext_ln823_174_fu_3814_p1 = $signed(p_Val2_875_fu_3804_p4);

assign sext_ln823_175_fu_9368_p1 = $signed(p_Val2_878_reg_11485);

assign sext_ln823_176_fu_9517_p1 = $signed(p_Val2_881_reg_11514);

assign sext_ln823_177_fu_9666_p1 = $signed(p_Val2_884_reg_11543);

assign sext_ln823_fu_2759_p1 = $signed(p_Val2_806_fu_2749_p4);

assign sext_ln856_153_fu_4107_p1 = p_Val2_810_reg_10812;

assign sext_ln856_154_fu_4353_p1 = p_Val2_816_reg_10874;

assign sext_ln856_155_fu_4478_p1 = p_Val2_819_reg_10905;

assign sext_ln856_156_fu_4603_p1 = p_Val2_822_reg_10936;

assign sext_ln856_157_fu_4728_p1 = p_Val2_825_reg_10967;

assign sext_ln856_158_fu_4853_p1 = p_Val2_828_reg_10998;

assign sext_ln856_159_fu_4978_p1 = p_Val2_831_reg_11029;

assign sext_ln856_160_fu_5115_p1 = p_Val2_834_fu_5109_p2;

assign sext_ln856_161_fu_5264_p1 = p_Val2_837_fu_5258_p2;

assign sext_ln856_162_fu_5413_p1 = p_Val2_840_fu_5407_p2;

assign sext_ln856_163_fu_5562_p1 = p_Val2_843_fu_5556_p2;

assign sext_ln856_164_fu_5711_p1 = p_Val2_846_fu_5705_p2;

assign sext_ln856_165_fu_5860_p1 = p_Val2_849_fu_5854_p2;

assign sext_ln856_166_fu_6009_p1 = p_Val2_852_fu_6003_p2;

assign sext_ln856_167_fu_6158_p1 = p_Val2_855_fu_6152_p2;

assign sext_ln856_168_fu_6307_p1 = p_Val2_858_fu_6301_p2;

assign sext_ln856_169_fu_8618_p1 = p_Val2_861_fu_8612_p2;

assign sext_ln856_170_fu_8767_p1 = p_Val2_864_fu_8761_p2;

assign sext_ln856_171_fu_8916_p1 = p_Val2_867_fu_8910_p2;

assign sext_ln856_172_fu_9065_p1 = p_Val2_870_fu_9059_p2;

assign sext_ln856_173_fu_9214_p1 = p_Val2_873_fu_9208_p2;

assign sext_ln856_174_fu_9351_p1 = p_Val2_876_reg_11319_pp0_iter1_reg;

assign sext_ln856_175_fu_9380_p1 = p_Val2_879_fu_9374_p2;

assign sext_ln856_176_fu_9529_p1 = p_Val2_882_fu_9523_p2;

assign sext_ln856_177_fu_9678_p1 = p_Val2_885_fu_9672_p2;

assign sext_ln856_fu_3982_p1 = p_Val2_807_reg_10781;

assign shl_ln_fu_3760_p3 = {{tmp288_fu_3750_p4}, {6'd0}};

assign tmp288_fu_3750_p4 = {{p_read_int_reg[95:64]}};

assign tmp_1287_fu_4010_p3 = r_V_178_reg_2283[32'd42];

assign tmp_1290_fu_2835_p3 = r_V_179_fu_262_p2[32'd23];

assign tmp_1293_fu_4135_p3 = r_V_179_reg_2287[32'd43];

assign tmp_1296_fu_2895_p3 = r_V_180_fu_251_p2[32'd23];

assign tmp_1299_fu_4257_p3 = r_V_180_reg_2291[32'd56];

assign tmp_1302_fu_2959_p3 = r_V_181_fu_256_p2[32'd23];

assign tmp_1305_fu_4381_p3 = r_V_181_reg_2295[32'd43];

assign tmp_1308_fu_3023_p3 = r_V_182_fu_264_p2[32'd23];

assign tmp_1311_fu_4506_p3 = r_V_182_reg_2299[32'd46];

assign tmp_1314_fu_3087_p3 = r_V_183_fu_240_p2[32'd23];

assign tmp_1317_fu_4631_p3 = r_V_183_reg_2303[32'd42];

assign tmp_1320_fu_3151_p3 = r_V_184_fu_249_p2[32'd23];

assign tmp_1323_fu_4756_p3 = r_V_184_reg_2307[32'd42];

assign tmp_1326_fu_3215_p3 = r_V_185_fu_259_p2[32'd23];

assign tmp_1329_fu_4881_p3 = r_V_185_reg_2311[32'd53];

assign tmp_1332_fu_3279_p3 = r_V_186_fu_246_p2[32'd23];

assign tmp_1335_fu_5006_p3 = r_V_186_reg_2315[32'd53];

assign tmp_1341_fu_5154_p3 = r_V_187_reg_2319[32'd40];

assign tmp_1347_fu_5303_p3 = r_V_188_reg_2323[32'd42];

assign tmp_1353_fu_5452_p3 = r_V_189_reg_2327[32'd44];

assign tmp_1359_fu_5601_p3 = r_V_190_reg_2331[32'd42];

assign tmp_1365_fu_5750_p3 = r_V_191_reg_2335[32'd53];

assign tmp_1371_fu_5899_p3 = r_V_192_reg_2339[32'd42];

assign tmp_1377_fu_6048_p3 = r_V_193_reg_2343[32'd42];

assign tmp_1383_fu_6197_p3 = r_V_194_reg_2347[32'd53];

assign tmp_1389_fu_6346_p3 = r_V_195_reg_2351[32'd53];

assign tmp_1395_fu_8657_p3 = r_V_reg_2675[32'd42];

assign tmp_1401_fu_8806_p3 = r_V_196_reg_2679[32'd41];

assign tmp_1407_fu_8955_p3 = r_V_197_reg_2683[32'd43];

assign tmp_1413_fu_9104_p3 = r_V_198_reg_2687[32'd44];

assign tmp_1419_fu_9253_p3 = r_V_199_reg_2691[32'd53];

assign tmp_1422_fu_3832_p3 = add_ln823_fu_3818_p2[32'd23];

assign tmp_1425_fu_3896_p3 = r_V_200_fu_3790_p2[32'd38];

assign tmp_1431_fu_9419_p3 = r_V_201_reg_2695[32'd40];

assign tmp_1437_fu_9568_p3 = r_V_202_reg_2699[32'd53];

assign tmp_1443_fu_9717_p3 = r_V_203_reg_2703[32'd53];

assign tmp_fu_2771_p3 = r_V_178_fu_254_p2[32'd23];

assign tmp_s_fu_3772_p4 = {{p_read_int_reg[81:64]}};

assign trunc_ln7_fu_3782_p3 = {{tmp_s_fu_3772_p4}, {6'd0}};

assign underflow_323_fu_4205_p2 = (xor_ln896_567_fu_4199_p2 & p_Result_809_reg_10800);

assign underflow_324_fu_4327_p2 = (xor_ln896_568_fu_4321_p2 & p_Result_812_reg_10831);

assign underflow_325_fu_4451_p2 = (xor_ln896_569_fu_4445_p2 & p_Result_815_reg_10862);

assign underflow_326_fu_4576_p2 = (xor_ln896_570_fu_4570_p2 & p_Result_818_reg_10893);

assign underflow_327_fu_4701_p2 = (xor_ln896_571_fu_4695_p2 & p_Result_821_reg_10924);

assign underflow_328_fu_4826_p2 = (xor_ln896_572_fu_4820_p2 & p_Result_824_reg_10955);

assign underflow_329_fu_4951_p2 = (xor_ln896_573_fu_4945_p2 & p_Result_827_reg_10986);

assign underflow_330_fu_5076_p2 = (xor_ln896_574_fu_5070_p2 & p_Result_830_reg_11017);

assign underflow_331_fu_5225_p2 = (xor_ln896_575_fu_5219_p2 & p_Result_833_reg_11048);

assign underflow_332_fu_5374_p2 = (xor_ln896_576_fu_5368_p2 & p_Result_836_reg_11077);

assign underflow_333_fu_5523_p2 = (xor_ln896_577_fu_5517_p2 & p_Result_839_reg_11106);

assign underflow_334_fu_5672_p2 = (xor_ln896_578_fu_5666_p2 & p_Result_842_reg_11135);

assign underflow_335_fu_5821_p2 = (xor_ln896_579_fu_5815_p2 & p_Result_845_reg_11164);

assign underflow_336_fu_5970_p2 = (xor_ln896_580_fu_5964_p2 & p_Result_848_reg_11193);

assign underflow_337_fu_6119_p2 = (xor_ln896_581_fu_6113_p2 & p_Result_851_reg_11222);

assign underflow_338_fu_6268_p2 = (xor_ln896_582_fu_6262_p2 & p_Result_854_reg_11251);

assign underflow_339_fu_6417_p2 = (xor_ln896_583_fu_6411_p2 & p_Result_857_reg_11280);

assign underflow_340_fu_8728_p2 = (xor_ln896_584_fu_8722_p2 & p_Result_860_reg_11334);

assign underflow_341_fu_8877_p2 = (xor_ln896_585_fu_8871_p2 & p_Result_863_reg_11363);

assign underflow_342_fu_9026_p2 = (xor_ln896_586_fu_9020_p2 & p_Result_866_reg_11392);

assign underflow_343_fu_9175_p2 = (xor_ln896_587_fu_9169_p2 & p_Result_869_reg_11421);

assign underflow_344_fu_9324_p2 = (xor_ln896_588_fu_9318_p2 & p_Result_872_reg_11450);

assign underflow_345_fu_3970_p2 = (xor_ln896_589_fu_3964_p2 & p_Result_875_fu_3796_p3);

assign underflow_346_fu_9490_p2 = (xor_ln896_590_fu_9484_p2 & p_Result_878_reg_11479);

assign underflow_347_fu_9639_p2 = (xor_ln896_591_fu_9633_p2 & p_Result_881_reg_11508);

assign underflow_348_fu_9788_p2 = (xor_ln896_592_fu_9782_p2 & p_Result_884_reg_11537);

assign underflow_349_fu_6856_p2 = (xor_ln896_538_fu_6850_p2 & p_Result_887_fu_6816_p3);

assign underflow_350_fu_6954_p2 = (xor_ln896_539_fu_6948_p2 & p_Result_889_fu_6914_p3);

assign underflow_351_fu_7052_p2 = (xor_ln896_540_fu_7046_p2 & p_Result_891_fu_7012_p3);

assign underflow_352_fu_7150_p2 = (xor_ln896_541_fu_7144_p2 & p_Result_893_fu_7110_p3);

assign underflow_353_fu_7248_p2 = (xor_ln896_542_fu_7242_p2 & p_Result_895_fu_7208_p3);

assign underflow_354_fu_7346_p2 = (xor_ln896_543_fu_7340_p2 & p_Result_897_fu_7306_p3);

assign underflow_355_fu_7444_p2 = (xor_ln896_544_fu_7438_p2 & p_Result_899_fu_7404_p3);

assign underflow_356_fu_7542_p2 = (xor_ln896_545_fu_7536_p2 & p_Result_901_fu_7502_p3);

assign underflow_357_fu_7640_p2 = (xor_ln896_546_fu_7634_p2 & p_Result_903_fu_7600_p3);

assign underflow_358_fu_7742_p2 = (xor_ln896_547_fu_7736_p2 & p_Result_905_fu_7702_p3);

assign underflow_359_fu_7844_p2 = (xor_ln896_548_fu_7838_p2 & p_Result_907_fu_7804_p3);

assign underflow_360_fu_7946_p2 = (xor_ln896_549_fu_7940_p2 & p_Result_909_fu_7906_p3);

assign underflow_361_fu_8048_p2 = (xor_ln896_550_fu_8042_p2 & p_Result_911_fu_8008_p3);

assign underflow_362_fu_8150_p2 = (xor_ln896_551_fu_8144_p2 & p_Result_913_fu_8110_p3);

assign underflow_363_fu_8252_p2 = (xor_ln896_552_fu_8246_p2 & p_Result_915_fu_8212_p3);

assign underflow_364_fu_8354_p2 = (xor_ln896_553_fu_8348_p2 & p_Result_917_fu_8314_p3);

assign underflow_365_fu_8456_p2 = (xor_ln896_554_fu_8450_p2 & p_Result_919_fu_8416_p3);

assign underflow_366_fu_8558_p2 = (xor_ln896_555_fu_8552_p2 & p_Result_921_fu_8518_p3);

assign underflow_367_fu_9867_p2 = (xor_ln896_556_fu_9861_p2 & p_Result_923_fu_9828_p3);

assign underflow_368_fu_9967_p2 = (xor_ln896_557_fu_9961_p2 & p_Result_925_fu_9928_p3);

assign underflow_369_fu_10067_p2 = (xor_ln896_558_fu_10061_p2 & p_Result_927_fu_10028_p3);

assign underflow_370_fu_10167_p2 = (xor_ln896_559_fu_10161_p2 & p_Result_929_fu_10128_p3);

assign underflow_371_fu_10267_p2 = (xor_ln896_560_fu_10261_p2 & p_Result_931_fu_10228_p3);

assign underflow_372_fu_10367_p2 = (xor_ln896_561_fu_10361_p2 & p_Result_933_fu_10328_p3);

assign underflow_373_fu_10467_p2 = (xor_ln896_562_fu_10461_p2 & p_Result_935_fu_10428_p3);

assign underflow_374_fu_10567_p2 = (xor_ln896_563_fu_10561_p2 & p_Result_937_fu_10528_p3);

assign underflow_375_fu_10667_p2 = (xor_ln896_564_fu_10661_p2 & p_Result_939_fu_10628_p3);

assign underflow_fu_4080_p2 = (xor_ln896_566_fu_4074_p2 & p_Result_s_reg_10769);

assign xor_ln302_323_fu_6868_p2 = (xor_ln302_fu_6862_p2 ^ 1'd1);

assign xor_ln302_324_fu_6960_p2 = (p_Result_890_fu_6928_p3 ^ p_Result_889_fu_6914_p3);

assign xor_ln302_325_fu_6966_p2 = (xor_ln302_324_fu_6960_p2 ^ 1'd1);

assign xor_ln302_326_fu_7058_p2 = (p_Result_892_fu_7026_p3 ^ p_Result_891_fu_7012_p3);

assign xor_ln302_327_fu_7064_p2 = (xor_ln302_326_fu_7058_p2 ^ 1'd1);

assign xor_ln302_328_fu_7156_p2 = (p_Result_894_fu_7124_p3 ^ p_Result_893_fu_7110_p3);

assign xor_ln302_329_fu_7162_p2 = (xor_ln302_328_fu_7156_p2 ^ 1'd1);

assign xor_ln302_330_fu_7254_p2 = (p_Result_896_fu_7222_p3 ^ p_Result_895_fu_7208_p3);

assign xor_ln302_331_fu_7260_p2 = (xor_ln302_330_fu_7254_p2 ^ 1'd1);

assign xor_ln302_332_fu_7352_p2 = (p_Result_898_fu_7320_p3 ^ p_Result_897_fu_7306_p3);

assign xor_ln302_333_fu_7358_p2 = (xor_ln302_332_fu_7352_p2 ^ 1'd1);

assign xor_ln302_334_fu_7450_p2 = (p_Result_900_fu_7418_p3 ^ p_Result_899_fu_7404_p3);

assign xor_ln302_335_fu_7456_p2 = (xor_ln302_334_fu_7450_p2 ^ 1'd1);

assign xor_ln302_336_fu_7548_p2 = (p_Result_902_fu_7516_p3 ^ p_Result_901_fu_7502_p3);

assign xor_ln302_337_fu_7554_p2 = (xor_ln302_336_fu_7548_p2 ^ 1'd1);

assign xor_ln302_338_fu_7646_p2 = (p_Result_904_fu_7614_p3 ^ p_Result_903_fu_7600_p3);

assign xor_ln302_339_fu_7652_p2 = (xor_ln302_338_fu_7646_p2 ^ 1'd1);

assign xor_ln302_340_fu_7748_p2 = (p_Result_906_fu_7716_p3 ^ p_Result_905_fu_7702_p3);

assign xor_ln302_341_fu_7754_p2 = (xor_ln302_340_fu_7748_p2 ^ 1'd1);

assign xor_ln302_342_fu_7850_p2 = (p_Result_908_fu_7818_p3 ^ p_Result_907_fu_7804_p3);

assign xor_ln302_343_fu_7856_p2 = (xor_ln302_342_fu_7850_p2 ^ 1'd1);

assign xor_ln302_344_fu_7952_p2 = (p_Result_910_fu_7920_p3 ^ p_Result_909_fu_7906_p3);

assign xor_ln302_345_fu_7958_p2 = (xor_ln302_344_fu_7952_p2 ^ 1'd1);

assign xor_ln302_346_fu_8054_p2 = (p_Result_912_fu_8022_p3 ^ p_Result_911_fu_8008_p3);

assign xor_ln302_347_fu_8060_p2 = (xor_ln302_346_fu_8054_p2 ^ 1'd1);

assign xor_ln302_348_fu_8156_p2 = (p_Result_914_fu_8124_p3 ^ p_Result_913_fu_8110_p3);

assign xor_ln302_349_fu_8162_p2 = (xor_ln302_348_fu_8156_p2 ^ 1'd1);

assign xor_ln302_350_fu_8258_p2 = (p_Result_916_fu_8226_p3 ^ p_Result_915_fu_8212_p3);

assign xor_ln302_351_fu_8264_p2 = (xor_ln302_350_fu_8258_p2 ^ 1'd1);

assign xor_ln302_352_fu_8360_p2 = (p_Result_918_fu_8328_p3 ^ p_Result_917_fu_8314_p3);

assign xor_ln302_353_fu_8366_p2 = (xor_ln302_352_fu_8360_p2 ^ 1'd1);

assign xor_ln302_354_fu_8462_p2 = (p_Result_920_fu_8430_p3 ^ p_Result_919_fu_8416_p3);

assign xor_ln302_355_fu_8468_p2 = (xor_ln302_354_fu_8462_p2 ^ 1'd1);

assign xor_ln302_356_fu_8564_p2 = (p_Result_922_fu_8532_p3 ^ p_Result_921_fu_8518_p3);

assign xor_ln302_357_fu_8570_p2 = (xor_ln302_356_fu_8564_p2 ^ 1'd1);

assign xor_ln302_358_fu_9873_p2 = (p_Result_924_fu_9841_p3 ^ p_Result_923_fu_9828_p3);

assign xor_ln302_359_fu_9879_p2 = (xor_ln302_358_fu_9873_p2 ^ 1'd1);

assign xor_ln302_360_fu_9973_p2 = (p_Result_926_fu_9941_p3 ^ p_Result_925_fu_9928_p3);

assign xor_ln302_361_fu_9979_p2 = (xor_ln302_360_fu_9973_p2 ^ 1'd1);

assign xor_ln302_362_fu_10073_p2 = (p_Result_928_fu_10041_p3 ^ p_Result_927_fu_10028_p3);

assign xor_ln302_363_fu_10079_p2 = (xor_ln302_362_fu_10073_p2 ^ 1'd1);

assign xor_ln302_364_fu_10173_p2 = (p_Result_930_fu_10141_p3 ^ p_Result_929_fu_10128_p3);

assign xor_ln302_365_fu_10179_p2 = (xor_ln302_364_fu_10173_p2 ^ 1'd1);

assign xor_ln302_366_fu_10273_p2 = (p_Result_932_fu_10241_p3 ^ p_Result_931_fu_10228_p3);

assign xor_ln302_367_fu_10279_p2 = (xor_ln302_366_fu_10273_p2 ^ 1'd1);

assign xor_ln302_368_fu_10373_p2 = (p_Result_934_fu_10341_p3 ^ p_Result_933_fu_10328_p3);

assign xor_ln302_369_fu_10379_p2 = (xor_ln302_368_fu_10373_p2 ^ 1'd1);

assign xor_ln302_370_fu_10473_p2 = (p_Result_936_fu_10441_p3 ^ p_Result_935_fu_10428_p3);

assign xor_ln302_371_fu_10479_p2 = (xor_ln302_370_fu_10473_p2 ^ 1'd1);

assign xor_ln302_372_fu_10573_p2 = (p_Result_938_fu_10541_p3 ^ p_Result_937_fu_10528_p3);

assign xor_ln302_373_fu_10579_p2 = (xor_ln302_372_fu_10573_p2 ^ 1'd1);

assign xor_ln302_374_fu_10673_p2 = (p_Result_940_fu_10641_p3 ^ p_Result_939_fu_10628_p3);

assign xor_ln302_375_fu_10679_p2 = (xor_ln302_374_fu_10673_p2 ^ 1'd1);

assign xor_ln302_fu_6862_p2 = (p_Result_888_fu_6830_p3 ^ p_Result_887_fu_6816_p3);

assign xor_ln888_321_fu_4120_p2 = (p_Result_810_reg_10806 ^ 1'd1);

assign xor_ln888_323_fu_4242_p2 = (p_Result_813_reg_10837 ^ 1'd1);

assign xor_ln888_325_fu_4366_p2 = (p_Result_816_reg_10868 ^ 1'd1);

assign xor_ln888_327_fu_4491_p2 = (p_Result_819_reg_10899 ^ 1'd1);

assign xor_ln888_329_fu_4616_p2 = (p_Result_822_reg_10930 ^ 1'd1);

assign xor_ln888_331_fu_4741_p2 = (p_Result_825_reg_10961 ^ 1'd1);

assign xor_ln888_333_fu_4866_p2 = (p_Result_828_reg_10992 ^ 1'd1);

assign xor_ln888_335_fu_4991_p2 = (p_Result_831_reg_11023 ^ 1'd1);

assign xor_ln888_337_fu_5138_p2 = (p_Result_834_reg_11059 ^ 1'd1);

assign xor_ln888_339_fu_5287_p2 = (p_Result_837_reg_11088 ^ 1'd1);

assign xor_ln888_341_fu_5436_p2 = (p_Result_840_reg_11117 ^ 1'd1);

assign xor_ln888_343_fu_5585_p2 = (p_Result_843_reg_11146 ^ 1'd1);

assign xor_ln888_345_fu_5734_p2 = (p_Result_846_reg_11175 ^ 1'd1);

assign xor_ln888_347_fu_5883_p2 = (p_Result_849_reg_11204 ^ 1'd1);

assign xor_ln888_349_fu_6032_p2 = (p_Result_852_reg_11233 ^ 1'd1);

assign xor_ln888_351_fu_6181_p2 = (p_Result_855_reg_11262 ^ 1'd1);

assign xor_ln888_353_fu_6330_p2 = (p_Result_858_reg_11291 ^ 1'd1);

assign xor_ln888_355_fu_8641_p2 = (p_Result_861_reg_11345 ^ 1'd1);

assign xor_ln888_357_fu_8790_p2 = (p_Result_864_reg_11374 ^ 1'd1);

assign xor_ln888_359_fu_8939_p2 = (p_Result_867_reg_11403 ^ 1'd1);

assign xor_ln888_361_fu_9088_p2 = (p_Result_870_reg_11432 ^ 1'd1);

assign xor_ln888_363_fu_9237_p2 = (p_Result_873_reg_11461 ^ 1'd1);

assign xor_ln888_365_fu_3878_p2 = (p_Result_876_fu_3824_p3 ^ 1'd1);

assign xor_ln888_367_fu_9403_p2 = (p_Result_879_reg_11490 ^ 1'd1);

assign xor_ln888_369_fu_9552_p2 = (p_Result_882_reg_11519 ^ 1'd1);

assign xor_ln888_371_fu_9701_p2 = (p_Result_885_reg_11548 ^ 1'd1);

assign xor_ln888_fu_3995_p2 = (p_Result_807_reg_10775 ^ 1'd1);

assign xor_ln890_159_fu_4143_p2 = (tmp_1293_fu_4135_p3 ^ 1'd1);

assign xor_ln890_160_fu_4265_p2 = (tmp_1299_fu_4257_p3 ^ 1'd1);

assign xor_ln890_161_fu_4389_p2 = (tmp_1305_fu_4381_p3 ^ 1'd1);

assign xor_ln890_162_fu_4514_p2 = (tmp_1311_fu_4506_p3 ^ 1'd1);

assign xor_ln890_163_fu_4639_p2 = (tmp_1317_fu_4631_p3 ^ 1'd1);

assign xor_ln890_164_fu_4764_p2 = (tmp_1323_fu_4756_p3 ^ 1'd1);

assign xor_ln890_165_fu_4889_p2 = (tmp_1329_fu_4881_p3 ^ 1'd1);

assign xor_ln890_166_fu_5014_p2 = (tmp_1335_fu_5006_p3 ^ 1'd1);

assign xor_ln890_167_fu_5162_p2 = (tmp_1341_fu_5154_p3 ^ 1'd1);

assign xor_ln890_168_fu_5311_p2 = (tmp_1347_fu_5303_p3 ^ 1'd1);

assign xor_ln890_169_fu_5460_p2 = (tmp_1353_fu_5452_p3 ^ 1'd1);

assign xor_ln890_170_fu_5609_p2 = (tmp_1359_fu_5601_p3 ^ 1'd1);

assign xor_ln890_171_fu_5758_p2 = (tmp_1365_fu_5750_p3 ^ 1'd1);

assign xor_ln890_172_fu_5907_p2 = (tmp_1371_fu_5899_p3 ^ 1'd1);

assign xor_ln890_173_fu_6056_p2 = (tmp_1377_fu_6048_p3 ^ 1'd1);

assign xor_ln890_174_fu_6205_p2 = (tmp_1383_fu_6197_p3 ^ 1'd1);

assign xor_ln890_175_fu_6354_p2 = (tmp_1389_fu_6346_p3 ^ 1'd1);

assign xor_ln890_176_fu_8665_p2 = (tmp_1395_fu_8657_p3 ^ 1'd1);

assign xor_ln890_177_fu_8814_p2 = (tmp_1401_fu_8806_p3 ^ 1'd1);

assign xor_ln890_178_fu_8963_p2 = (tmp_1407_fu_8955_p3 ^ 1'd1);

assign xor_ln890_179_fu_9112_p2 = (tmp_1413_fu_9104_p3 ^ 1'd1);

assign xor_ln890_180_fu_9261_p2 = (tmp_1419_fu_9253_p3 ^ 1'd1);

assign xor_ln890_181_fu_3904_p2 = (tmp_1425_fu_3896_p3 ^ 1'd1);

assign xor_ln890_182_fu_9427_p2 = (tmp_1431_fu_9419_p3 ^ 1'd1);

assign xor_ln890_183_fu_9576_p2 = (tmp_1437_fu_9568_p3 ^ 1'd1);

assign xor_ln890_184_fu_9725_p2 = (tmp_1443_fu_9717_p3 ^ 1'd1);

assign xor_ln890_fu_4018_p2 = (tmp_1287_fu_4010_p3 ^ 1'd1);

assign xor_ln895_485_fu_4051_p2 = (p_Result_s_reg_10769 ^ 1'd1);

assign xor_ln895_486_fu_4165_p2 = (deleted_zeros_158_fu_4130_p2 ^ 1'd1);

assign xor_ln895_487_fu_4176_p2 = (p_Result_809_reg_10800 ^ 1'd1);

assign xor_ln895_488_fu_4287_p2 = (deleted_zeros_159_fu_4252_p2 ^ 1'd1);

assign xor_ln895_489_fu_4298_p2 = (p_Result_812_reg_10831 ^ 1'd1);

assign xor_ln895_490_fu_4411_p2 = (deleted_zeros_160_fu_4376_p2 ^ 1'd1);

assign xor_ln895_491_fu_4422_p2 = (p_Result_815_reg_10862 ^ 1'd1);

assign xor_ln895_492_fu_4536_p2 = (deleted_zeros_161_fu_4501_p2 ^ 1'd1);

assign xor_ln895_493_fu_4547_p2 = (p_Result_818_reg_10893 ^ 1'd1);

assign xor_ln895_494_fu_4661_p2 = (deleted_zeros_162_fu_4626_p2 ^ 1'd1);

assign xor_ln895_495_fu_4672_p2 = (p_Result_821_reg_10924 ^ 1'd1);

assign xor_ln895_496_fu_4786_p2 = (deleted_zeros_163_fu_4751_p2 ^ 1'd1);

assign xor_ln895_497_fu_4797_p2 = (p_Result_824_reg_10955 ^ 1'd1);

assign xor_ln895_498_fu_4911_p2 = (deleted_zeros_164_fu_4876_p2 ^ 1'd1);

assign xor_ln895_499_fu_4922_p2 = (p_Result_827_reg_10986 ^ 1'd1);

assign xor_ln895_500_fu_5036_p2 = (deleted_zeros_165_fu_5001_p2 ^ 1'd1);

assign xor_ln895_501_fu_5047_p2 = (p_Result_830_reg_11017 ^ 1'd1);

assign xor_ln895_502_fu_5184_p2 = (deleted_zeros_166_fu_5149_p2 ^ 1'd1);

assign xor_ln895_503_fu_5196_p2 = (p_Result_833_reg_11048 ^ 1'd1);

assign xor_ln895_504_fu_5333_p2 = (deleted_zeros_167_fu_5298_p2 ^ 1'd1);

assign xor_ln895_505_fu_5345_p2 = (p_Result_836_reg_11077 ^ 1'd1);

assign xor_ln895_506_fu_5482_p2 = (deleted_zeros_168_fu_5447_p2 ^ 1'd1);

assign xor_ln895_507_fu_5494_p2 = (p_Result_839_reg_11106 ^ 1'd1);

assign xor_ln895_508_fu_5631_p2 = (deleted_zeros_169_fu_5596_p2 ^ 1'd1);

assign xor_ln895_509_fu_5643_p2 = (p_Result_842_reg_11135 ^ 1'd1);

assign xor_ln895_510_fu_5780_p2 = (deleted_zeros_170_fu_5745_p2 ^ 1'd1);

assign xor_ln895_511_fu_5792_p2 = (p_Result_845_reg_11164 ^ 1'd1);

assign xor_ln895_512_fu_5929_p2 = (deleted_zeros_171_fu_5894_p2 ^ 1'd1);

assign xor_ln895_513_fu_5941_p2 = (p_Result_848_reg_11193 ^ 1'd1);

assign xor_ln895_514_fu_6078_p2 = (deleted_zeros_172_fu_6043_p2 ^ 1'd1);

assign xor_ln895_515_fu_6090_p2 = (p_Result_851_reg_11222 ^ 1'd1);

assign xor_ln895_516_fu_6227_p2 = (deleted_zeros_173_fu_6192_p2 ^ 1'd1);

assign xor_ln895_517_fu_6239_p2 = (p_Result_854_reg_11251 ^ 1'd1);

assign xor_ln895_518_fu_6376_p2 = (deleted_zeros_174_fu_6341_p2 ^ 1'd1);

assign xor_ln895_519_fu_6388_p2 = (p_Result_857_reg_11280 ^ 1'd1);

assign xor_ln895_520_fu_8687_p2 = (deleted_zeros_175_fu_8652_p2 ^ 1'd1);

assign xor_ln895_521_fu_8699_p2 = (p_Result_860_reg_11334 ^ 1'd1);

assign xor_ln895_522_fu_8836_p2 = (deleted_zeros_176_fu_8801_p2 ^ 1'd1);

assign xor_ln895_523_fu_8848_p2 = (p_Result_863_reg_11363 ^ 1'd1);

assign xor_ln895_524_fu_8985_p2 = (deleted_zeros_177_fu_8950_p2 ^ 1'd1);

assign xor_ln895_525_fu_8997_p2 = (p_Result_866_reg_11392 ^ 1'd1);

assign xor_ln895_526_fu_9134_p2 = (deleted_zeros_178_fu_9099_p2 ^ 1'd1);

assign xor_ln895_527_fu_9146_p2 = (p_Result_869_reg_11421 ^ 1'd1);

assign xor_ln895_528_fu_9283_p2 = (deleted_zeros_179_fu_9248_p2 ^ 1'd1);

assign xor_ln895_529_fu_9295_p2 = (p_Result_872_reg_11450 ^ 1'd1);

assign xor_ln895_530_fu_3928_p2 = (deleted_zeros_180_fu_3890_p2 ^ 1'd1);

assign xor_ln895_531_fu_3940_p2 = (p_Result_875_fu_3796_p3 ^ 1'd1);

assign xor_ln895_532_fu_9449_p2 = (deleted_zeros_181_fu_9414_p2 ^ 1'd1);

assign xor_ln895_533_fu_9461_p2 = (p_Result_878_reg_11479 ^ 1'd1);

assign xor_ln895_534_fu_9598_p2 = (deleted_zeros_182_fu_9563_p2 ^ 1'd1);

assign xor_ln895_535_fu_9610_p2 = (p_Result_881_reg_11508 ^ 1'd1);

assign xor_ln895_536_fu_9747_p2 = (deleted_zeros_183_fu_9712_p2 ^ 1'd1);

assign xor_ln895_537_fu_9759_p2 = (p_Result_884_reg_11537 ^ 1'd1);

assign xor_ln895_538_fu_6838_p2 = (p_Result_887_fu_6816_p3 ^ 1'd1);

assign xor_ln895_539_fu_6936_p2 = (p_Result_889_fu_6914_p3 ^ 1'd1);

assign xor_ln895_540_fu_7034_p2 = (p_Result_891_fu_7012_p3 ^ 1'd1);

assign xor_ln895_541_fu_7132_p2 = (p_Result_893_fu_7110_p3 ^ 1'd1);

assign xor_ln895_542_fu_7230_p2 = (p_Result_895_fu_7208_p3 ^ 1'd1);

assign xor_ln895_543_fu_7328_p2 = (p_Result_897_fu_7306_p3 ^ 1'd1);

assign xor_ln895_544_fu_7426_p2 = (p_Result_899_fu_7404_p3 ^ 1'd1);

assign xor_ln895_545_fu_7524_p2 = (p_Result_901_fu_7502_p3 ^ 1'd1);

assign xor_ln895_546_fu_7622_p2 = (p_Result_903_fu_7600_p3 ^ 1'd1);

assign xor_ln895_547_fu_7724_p2 = (p_Result_905_fu_7702_p3 ^ 1'd1);

assign xor_ln895_548_fu_7826_p2 = (p_Result_907_fu_7804_p3 ^ 1'd1);

assign xor_ln895_549_fu_7928_p2 = (p_Result_909_fu_7906_p3 ^ 1'd1);

assign xor_ln895_550_fu_8030_p2 = (p_Result_911_fu_8008_p3 ^ 1'd1);

assign xor_ln895_551_fu_8132_p2 = (p_Result_913_fu_8110_p3 ^ 1'd1);

assign xor_ln895_552_fu_8234_p2 = (p_Result_915_fu_8212_p3 ^ 1'd1);

assign xor_ln895_553_fu_8336_p2 = (p_Result_917_fu_8314_p3 ^ 1'd1);

assign xor_ln895_554_fu_8438_p2 = (p_Result_919_fu_8416_p3 ^ 1'd1);

assign xor_ln895_555_fu_8540_p2 = (p_Result_921_fu_8518_p3 ^ 1'd1);

assign xor_ln895_556_fu_9849_p2 = (p_Result_923_fu_9828_p3 ^ 1'd1);

assign xor_ln895_557_fu_9949_p2 = (p_Result_925_fu_9928_p3 ^ 1'd1);

assign xor_ln895_558_fu_10049_p2 = (p_Result_927_fu_10028_p3 ^ 1'd1);

assign xor_ln895_559_fu_10149_p2 = (p_Result_929_fu_10128_p3 ^ 1'd1);

assign xor_ln895_560_fu_10249_p2 = (p_Result_931_fu_10228_p3 ^ 1'd1);

assign xor_ln895_561_fu_10349_p2 = (p_Result_933_fu_10328_p3 ^ 1'd1);

assign xor_ln895_562_fu_10449_p2 = (p_Result_935_fu_10428_p3 ^ 1'd1);

assign xor_ln895_563_fu_10549_p2 = (p_Result_937_fu_10528_p3 ^ 1'd1);

assign xor_ln895_564_fu_10649_p2 = (p_Result_939_fu_10628_p3 ^ 1'd1);

assign xor_ln895_fu_4040_p2 = (deleted_zeros_fu_4005_p2 ^ 1'd1);

assign xor_ln896_485_fu_4062_p2 = (deleted_ones_fu_4030_p2 ^ 1'd1);

assign xor_ln896_486_fu_4110_p2 = (p_Result_811_reg_10817 ^ 1'd1);

assign xor_ln896_487_fu_4187_p2 = (deleted_ones_323_fu_4155_p2 ^ 1'd1);

assign xor_ln896_488_fu_4232_p2 = (p_Result_814_reg_10848 ^ 1'd1);

assign xor_ln896_489_fu_4309_p2 = (deleted_ones_324_fu_4277_p2 ^ 1'd1);

assign xor_ln896_490_fu_4356_p2 = (p_Result_817_reg_10879 ^ 1'd1);

assign xor_ln896_491_fu_4433_p2 = (deleted_ones_325_fu_4401_p2 ^ 1'd1);

assign xor_ln896_492_fu_4481_p2 = (p_Result_820_reg_10910 ^ 1'd1);

assign xor_ln896_493_fu_4558_p2 = (deleted_ones_326_fu_4526_p2 ^ 1'd1);

assign xor_ln896_494_fu_4606_p2 = (p_Result_823_reg_10941 ^ 1'd1);

assign xor_ln896_495_fu_4683_p2 = (deleted_ones_327_fu_4651_p2 ^ 1'd1);

assign xor_ln896_496_fu_4731_p2 = (p_Result_826_reg_10972 ^ 1'd1);

assign xor_ln896_497_fu_4808_p2 = (deleted_ones_328_fu_4776_p2 ^ 1'd1);

assign xor_ln896_498_fu_4856_p2 = (p_Result_829_reg_11003 ^ 1'd1);

assign xor_ln896_499_fu_4933_p2 = (deleted_ones_329_fu_4901_p2 ^ 1'd1);

assign xor_ln896_500_fu_4981_p2 = (p_Result_832_reg_11034 ^ 1'd1);

assign xor_ln896_501_fu_5058_p2 = (deleted_ones_330_fu_5026_p2 ^ 1'd1);

assign xor_ln896_502_fu_5127_p2 = (p_Result_835_fu_5119_p3 ^ 1'd1);

assign xor_ln896_503_fu_5207_p2 = (deleted_ones_331_fu_5174_p2 ^ 1'd1);

assign xor_ln896_504_fu_5276_p2 = (p_Result_838_fu_5268_p3 ^ 1'd1);

assign xor_ln896_505_fu_5356_p2 = (deleted_ones_332_fu_5323_p2 ^ 1'd1);

assign xor_ln896_506_fu_5425_p2 = (p_Result_841_fu_5417_p3 ^ 1'd1);

assign xor_ln896_507_fu_5505_p2 = (deleted_ones_333_fu_5472_p2 ^ 1'd1);

assign xor_ln896_508_fu_5574_p2 = (p_Result_844_fu_5566_p3 ^ 1'd1);

assign xor_ln896_509_fu_5654_p2 = (deleted_ones_334_fu_5621_p2 ^ 1'd1);

assign xor_ln896_510_fu_5723_p2 = (p_Result_847_fu_5715_p3 ^ 1'd1);

assign xor_ln896_511_fu_5803_p2 = (deleted_ones_335_fu_5770_p2 ^ 1'd1);

assign xor_ln896_512_fu_5872_p2 = (p_Result_850_fu_5864_p3 ^ 1'd1);

assign xor_ln896_513_fu_5952_p2 = (deleted_ones_336_fu_5919_p2 ^ 1'd1);

assign xor_ln896_514_fu_6021_p2 = (p_Result_853_fu_6013_p3 ^ 1'd1);

assign xor_ln896_515_fu_6101_p2 = (deleted_ones_337_fu_6068_p2 ^ 1'd1);

assign xor_ln896_516_fu_6170_p2 = (p_Result_856_fu_6162_p3 ^ 1'd1);

assign xor_ln896_517_fu_6250_p2 = (deleted_ones_338_fu_6217_p2 ^ 1'd1);

assign xor_ln896_518_fu_6319_p2 = (p_Result_859_fu_6311_p3 ^ 1'd1);

assign xor_ln896_519_fu_6399_p2 = (deleted_ones_339_fu_6366_p2 ^ 1'd1);

assign xor_ln896_520_fu_8630_p2 = (p_Result_862_fu_8622_p3 ^ 1'd1);

assign xor_ln896_521_fu_8710_p2 = (deleted_ones_340_fu_8677_p2 ^ 1'd1);

assign xor_ln896_522_fu_8779_p2 = (p_Result_865_fu_8771_p3 ^ 1'd1);

assign xor_ln896_523_fu_8859_p2 = (deleted_ones_341_fu_8826_p2 ^ 1'd1);

assign xor_ln896_524_fu_8928_p2 = (p_Result_868_fu_8920_p3 ^ 1'd1);

assign xor_ln896_525_fu_9008_p2 = (deleted_ones_342_fu_8975_p2 ^ 1'd1);

assign xor_ln896_526_fu_9077_p2 = (p_Result_871_fu_9069_p3 ^ 1'd1);

assign xor_ln896_527_fu_9157_p2 = (deleted_ones_343_fu_9124_p2 ^ 1'd1);

assign xor_ln896_528_fu_9226_p2 = (p_Result_874_fu_9218_p3 ^ 1'd1);

assign xor_ln896_529_fu_9306_p2 = (deleted_ones_344_fu_9273_p2 ^ 1'd1);

assign xor_ln896_530_fu_3858_p2 = (p_Result_877_fu_3850_p3 ^ 1'd1);

assign xor_ln896_531_fu_3952_p2 = (deleted_ones_345_fu_3916_p2 ^ 1'd1);

assign xor_ln896_532_fu_9392_p2 = (p_Result_880_fu_9384_p3 ^ 1'd1);

assign xor_ln896_533_fu_9472_p2 = (deleted_ones_346_fu_9439_p2 ^ 1'd1);

assign xor_ln896_534_fu_9541_p2 = (p_Result_883_fu_9533_p3 ^ 1'd1);

assign xor_ln896_535_fu_9621_p2 = (deleted_ones_347_fu_9588_p2 ^ 1'd1);

assign xor_ln896_536_fu_9690_p2 = (p_Result_886_fu_9682_p3 ^ 1'd1);

assign xor_ln896_537_fu_9770_p2 = (deleted_ones_348_fu_9737_p2 ^ 1'd1);

assign xor_ln896_538_fu_6850_p2 = (p_Result_888_fu_6830_p3 ^ 1'd1);

assign xor_ln896_539_fu_6948_p2 = (p_Result_890_fu_6928_p3 ^ 1'd1);

assign xor_ln896_540_fu_7046_p2 = (p_Result_892_fu_7026_p3 ^ 1'd1);

assign xor_ln896_541_fu_7144_p2 = (p_Result_894_fu_7124_p3 ^ 1'd1);

assign xor_ln896_542_fu_7242_p2 = (p_Result_896_fu_7222_p3 ^ 1'd1);

assign xor_ln896_543_fu_7340_p2 = (p_Result_898_fu_7320_p3 ^ 1'd1);

assign xor_ln896_544_fu_7438_p2 = (p_Result_900_fu_7418_p3 ^ 1'd1);

assign xor_ln896_545_fu_7536_p2 = (p_Result_902_fu_7516_p3 ^ 1'd1);

assign xor_ln896_546_fu_7634_p2 = (p_Result_904_fu_7614_p3 ^ 1'd1);

assign xor_ln896_547_fu_7736_p2 = (p_Result_906_fu_7716_p3 ^ 1'd1);

assign xor_ln896_548_fu_7838_p2 = (p_Result_908_fu_7818_p3 ^ 1'd1);

assign xor_ln896_549_fu_7940_p2 = (p_Result_910_fu_7920_p3 ^ 1'd1);

assign xor_ln896_550_fu_8042_p2 = (p_Result_912_fu_8022_p3 ^ 1'd1);

assign xor_ln896_551_fu_8144_p2 = (p_Result_914_fu_8124_p3 ^ 1'd1);

assign xor_ln896_552_fu_8246_p2 = (p_Result_916_fu_8226_p3 ^ 1'd1);

assign xor_ln896_553_fu_8348_p2 = (p_Result_918_fu_8328_p3 ^ 1'd1);

assign xor_ln896_554_fu_8450_p2 = (p_Result_920_fu_8430_p3 ^ 1'd1);

assign xor_ln896_555_fu_8552_p2 = (p_Result_922_fu_8532_p3 ^ 1'd1);

assign xor_ln896_556_fu_9861_p2 = (p_Result_924_fu_9841_p3 ^ 1'd1);

assign xor_ln896_557_fu_9961_p2 = (p_Result_926_fu_9941_p3 ^ 1'd1);

assign xor_ln896_558_fu_10061_p2 = (p_Result_928_fu_10041_p3 ^ 1'd1);

assign xor_ln896_559_fu_10161_p2 = (p_Result_930_fu_10141_p3 ^ 1'd1);

assign xor_ln896_560_fu_10261_p2 = (p_Result_932_fu_10241_p3 ^ 1'd1);

assign xor_ln896_561_fu_10361_p2 = (p_Result_934_fu_10341_p3 ^ 1'd1);

assign xor_ln896_562_fu_10461_p2 = (p_Result_936_fu_10441_p3 ^ 1'd1);

assign xor_ln896_563_fu_10561_p2 = (p_Result_938_fu_10541_p3 ^ 1'd1);

assign xor_ln896_564_fu_10661_p2 = (p_Result_940_fu_10641_p3 ^ 1'd1);

assign xor_ln896_566_fu_4074_p2 = (or_ln896_fu_4068_p2 ^ and_ln891_fu_4035_p2);

assign xor_ln896_567_fu_4199_p2 = (or_ln896_161_fu_4193_p2 ^ and_ln891_161_fu_4160_p2);

assign xor_ln896_568_fu_4321_p2 = (or_ln896_162_fu_4315_p2 ^ and_ln891_162_fu_4282_p2);

assign xor_ln896_569_fu_4445_p2 = (or_ln896_163_fu_4439_p2 ^ and_ln891_163_fu_4406_p2);

assign xor_ln896_570_fu_4570_p2 = (or_ln896_164_fu_4564_p2 ^ and_ln891_164_fu_4531_p2);

assign xor_ln896_571_fu_4695_p2 = (or_ln896_165_fu_4689_p2 ^ and_ln891_165_fu_4656_p2);

assign xor_ln896_572_fu_4820_p2 = (or_ln896_166_fu_4814_p2 ^ and_ln891_166_fu_4781_p2);

assign xor_ln896_573_fu_4945_p2 = (or_ln896_167_fu_4939_p2 ^ and_ln891_167_fu_4906_p2);

assign xor_ln896_574_fu_5070_p2 = (or_ln896_168_fu_5064_p2 ^ and_ln891_168_fu_5031_p2);

assign xor_ln896_575_fu_5219_p2 = (or_ln896_169_fu_5213_p2 ^ and_ln891_169_fu_5179_p2);

assign xor_ln896_576_fu_5368_p2 = (or_ln896_170_fu_5362_p2 ^ and_ln891_170_fu_5328_p2);

assign xor_ln896_577_fu_5517_p2 = (or_ln896_171_fu_5511_p2 ^ and_ln891_171_fu_5477_p2);

assign xor_ln896_578_fu_5666_p2 = (or_ln896_172_fu_5660_p2 ^ and_ln891_172_fu_5626_p2);

assign xor_ln896_579_fu_5815_p2 = (or_ln896_173_fu_5809_p2 ^ and_ln891_173_fu_5775_p2);

assign xor_ln896_580_fu_5964_p2 = (or_ln896_174_fu_5958_p2 ^ and_ln891_174_fu_5924_p2);

assign xor_ln896_581_fu_6113_p2 = (or_ln896_175_fu_6107_p2 ^ and_ln891_175_fu_6073_p2);

assign xor_ln896_582_fu_6262_p2 = (or_ln896_176_fu_6256_p2 ^ and_ln891_176_fu_6222_p2);

assign xor_ln896_583_fu_6411_p2 = (or_ln896_177_fu_6405_p2 ^ and_ln891_177_fu_6371_p2);

assign xor_ln896_584_fu_8722_p2 = (or_ln896_178_fu_8716_p2 ^ and_ln891_178_fu_8682_p2);

assign xor_ln896_585_fu_8871_p2 = (or_ln896_179_fu_8865_p2 ^ and_ln891_179_fu_8831_p2);

assign xor_ln896_586_fu_9020_p2 = (or_ln896_180_fu_9014_p2 ^ and_ln891_180_fu_8980_p2);

assign xor_ln896_587_fu_9169_p2 = (or_ln896_181_fu_9163_p2 ^ and_ln891_181_fu_9129_p2);

assign xor_ln896_588_fu_9318_p2 = (or_ln896_182_fu_9312_p2 ^ and_ln891_182_fu_9278_p2);

assign xor_ln896_589_fu_3964_p2 = (or_ln896_183_fu_3958_p2 ^ and_ln891_183_fu_3922_p2);

assign xor_ln896_590_fu_9484_p2 = (or_ln896_184_fu_9478_p2 ^ and_ln891_184_fu_9444_p2);

assign xor_ln896_591_fu_9633_p2 = (or_ln896_185_fu_9627_p2 ^ and_ln891_185_fu_9593_p2);

assign xor_ln896_592_fu_9782_p2 = (or_ln896_186_fu_9776_p2 ^ and_ln891_186_fu_9742_p2);

assign xor_ln896_fu_3985_p2 = (p_Result_808_reg_10786 ^ 1'd1);

assign zext_ln377_161_fu_2843_p1 = tmp_1290_fu_2835_p3;

assign zext_ln377_162_fu_2903_p1 = tmp_1296_fu_2895_p3;

assign zext_ln377_163_fu_2967_p1 = tmp_1302_fu_2959_p3;

assign zext_ln377_164_fu_3031_p1 = tmp_1308_fu_3023_p3;

assign zext_ln377_165_fu_3095_p1 = tmp_1314_fu_3087_p3;

assign zext_ln377_166_fu_3159_p1 = tmp_1320_fu_3151_p3;

assign zext_ln377_167_fu_3223_p1 = tmp_1326_fu_3215_p3;

assign zext_ln377_168_fu_3287_p1 = tmp_1332_fu_3279_p3;

assign zext_ln377_169_fu_5106_p1 = tmp_1338_reg_11065;

assign zext_ln377_170_fu_5255_p1 = tmp_1344_reg_11094;

assign zext_ln377_171_fu_5404_p1 = tmp_1350_reg_11123;

assign zext_ln377_172_fu_5553_p1 = tmp_1356_reg_11152;

assign zext_ln377_173_fu_5702_p1 = tmp_1362_reg_11181;

assign zext_ln377_174_fu_5851_p1 = tmp_1368_reg_11210;

assign zext_ln377_175_fu_6000_p1 = tmp_1374_reg_11239;

assign zext_ln377_176_fu_6149_p1 = tmp_1380_reg_11268;

assign zext_ln377_177_fu_6298_p1 = tmp_1386_reg_11297;

assign zext_ln377_178_fu_8609_p1 = tmp_1392_reg_11351;

assign zext_ln377_179_fu_8758_p1 = tmp_1398_reg_11380;

assign zext_ln377_180_fu_8907_p1 = tmp_1404_reg_11409;

assign zext_ln377_181_fu_9056_p1 = tmp_1410_reg_11438;

assign zext_ln377_182_fu_9205_p1 = tmp_1416_reg_11467;

assign zext_ln377_183_fu_3840_p1 = tmp_1422_fu_3832_p3;

assign zext_ln377_184_fu_9371_p1 = tmp_1428_reg_11496;

assign zext_ln377_185_fu_9520_p1 = tmp_1434_reg_11525;

assign zext_ln377_186_fu_9669_p1 = tmp_1440_reg_11554;

assign zext_ln377_fu_2779_p1 = tmp_fu_2771_p3;

endmodule //motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config2_s
