module mpc_qp_admm_Pipeline_mvmult_row (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        temp1_V_3_04,
        temp1_V_2_03,
        temp1_V_1_02,
        temp1_V_0_01,
        sext_ln1273,
        sext_ln1273_1,
        sext_ln1273_24,
        sext_ln1273_3,
        sext_ln1273_4,
        sext_ln1273_5,
        sext_ln1273_6,
        sext_ln1273_7,
        sext_ln1273_8,
        sext_ln1273_9,
        sext_ln1273_10,
        sext_ln1273_11,
        sext_ln1273_12,
        sext_ln1273_13,
        sext_ln1273_14,
        sext_ln1273_15,
        sext_ln1273_16,
        sext_ln1273_17,
        sext_ln1273_18,
        sext_ln1273_19,
        sext_ln1273_20,
        sext_ln1273_21,
        sext_ln1273_22,
        sext_ln1273_23,
        temp1_V_3_1_out,
        temp1_V_3_1_out_ap_vld,
        temp1_V_2_1_out,
        temp1_V_2_1_out_ap_vld,
        temp1_V_1_1_out,
        temp1_V_1_1_out_ap_vld,
        temp1_V_0_1_out,
        temp1_V_0_1_out_ap_vld
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] temp1_V_3_04;
input  [31:0] temp1_V_2_03;
input  [31:0] temp1_V_1_02;
input  [31:0] temp1_V_0_01;
input  [31:0] sext_ln1273;
input  [31:0] sext_ln1273_1;
input  [31:0] sext_ln1273_24;
input  [31:0] sext_ln1273_3;
input  [31:0] sext_ln1273_4;
input  [31:0] sext_ln1273_5;
input  [31:0] sext_ln1273_6;
input  [31:0] sext_ln1273_7;
input  [31:0] sext_ln1273_8;
input  [31:0] sext_ln1273_9;
input  [31:0] sext_ln1273_10;
input  [31:0] sext_ln1273_11;
input  [31:0] sext_ln1273_12;
input  [31:0] sext_ln1273_13;
input  [31:0] sext_ln1273_14;
input  [31:0] sext_ln1273_15;
input  [31:0] sext_ln1273_16;
input  [31:0] sext_ln1273_17;
input  [31:0] sext_ln1273_18;
input  [31:0] sext_ln1273_19;
input  [31:0] sext_ln1273_20;
input  [31:0] sext_ln1273_21;
input  [31:0] sext_ln1273_22;
input  [31:0] sext_ln1273_23;
output  [31:0] temp1_V_3_1_out;
output   temp1_V_3_1_out_ap_vld;
output  [31:0] temp1_V_2_1_out;
output   temp1_V_2_1_out_ap_vld;
output  [31:0] temp1_V_1_1_out;
output   temp1_V_1_1_out_ap_vld;
output  [31:0] temp1_V_0_1_out;
output   temp1_V_0_1_out_ap_vld;

reg ap_idle;
reg temp1_V_3_1_out_ap_vld;
reg temp1_V_2_1_out_ap_vld;
reg temp1_V_1_1_out_ap_vld;
reg temp1_V_0_1_out_ap_vld;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
reg    ap_enable_reg_pp0_iter23;
reg    ap_enable_reg_pp0_iter24;
reg    ap_enable_reg_pp0_iter25;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_state21_pp0_stage0_iter20;
wire    ap_block_state22_pp0_stage0_iter21;
wire    ap_block_state23_pp0_stage0_iter22;
wire    ap_block_state24_pp0_stage0_iter23;
wire    ap_block_state25_pp0_stage0_iter24;
wire    ap_block_state26_pp0_stage0_iter25;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] icmp_ln24_fu_514_p2;
reg    ap_condition_exit_pp0_iter0_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire    ap_block_pp0_stage0_11001;
wire  signed [63:0] sext_ln1273_23_cast_fu_390_p1;
reg  signed [63:0] sext_ln1273_23_cast_reg_6498;
wire  signed [63:0] sext_ln1273_22_cast_fu_394_p1;
reg  signed [63:0] sext_ln1273_22_cast_reg_6503;
wire  signed [63:0] sext_ln1273_21_cast_fu_398_p1;
reg  signed [63:0] sext_ln1273_21_cast_reg_6508;
wire  signed [63:0] sext_ln1273_20_cast_fu_402_p1;
reg  signed [63:0] sext_ln1273_20_cast_reg_6513;
wire  signed [63:0] sext_ln1273_19_cast_fu_406_p1;
reg  signed [63:0] sext_ln1273_19_cast_reg_6518;
wire  signed [63:0] sext_ln1273_18_cast_fu_410_p1;
reg  signed [63:0] sext_ln1273_18_cast_reg_6523;
wire  signed [63:0] sext_ln1273_17_cast_fu_414_p1;
reg  signed [63:0] sext_ln1273_17_cast_reg_6528;
wire  signed [63:0] sext_ln1273_16_cast_fu_418_p1;
reg  signed [63:0] sext_ln1273_16_cast_reg_6533;
wire  signed [63:0] sext_ln1273_15_cast_fu_422_p1;
reg  signed [63:0] sext_ln1273_15_cast_reg_6538;
wire  signed [63:0] sext_ln1273_14_cast_fu_426_p1;
reg  signed [63:0] sext_ln1273_14_cast_reg_6543;
wire  signed [63:0] sext_ln1273_13_cast_fu_430_p1;
reg  signed [63:0] sext_ln1273_13_cast_reg_6548;
wire  signed [63:0] sext_ln1273_12_cast_fu_434_p1;
reg  signed [63:0] sext_ln1273_12_cast_reg_6553;
wire  signed [63:0] sext_ln1273_11_cast_fu_438_p1;
reg  signed [63:0] sext_ln1273_11_cast_reg_6558;
wire  signed [63:0] sext_ln1273_10_cast_fu_442_p1;
reg  signed [63:0] sext_ln1273_10_cast_reg_6563;
wire  signed [63:0] sext_ln1273_9_cast_fu_446_p1;
reg  signed [63:0] sext_ln1273_9_cast_reg_6568;
wire  signed [63:0] sext_ln1273_8_cast_fu_450_p1;
reg  signed [63:0] sext_ln1273_8_cast_reg_6573;
wire  signed [63:0] sext_ln1273_7_cast_fu_454_p1;
reg  signed [63:0] sext_ln1273_7_cast_reg_6578;
wire  signed [63:0] sext_ln1273_6_cast_fu_458_p1;
reg  signed [63:0] sext_ln1273_6_cast_reg_6583;
wire  signed [63:0] sext_ln1273_5_cast_fu_462_p1;
reg  signed [63:0] sext_ln1273_5_cast_reg_6588;
wire  signed [63:0] sext_ln1273_4_cast_fu_466_p1;
reg  signed [63:0] sext_ln1273_4_cast_reg_6593;
wire  signed [63:0] sext_ln1273_3_cast_fu_470_p1;
reg  signed [63:0] sext_ln1273_3_cast_reg_6598;
wire  signed [63:0] sext_ln1273_24_cast_fu_474_p1;
reg  signed [63:0] sext_ln1273_24_cast_reg_6603;
wire  signed [63:0] sext_ln1273_1_cast_fu_478_p1;
reg  signed [63:0] sext_ln1273_1_cast_reg_6608;
wire  signed [63:0] sext_ln1273_cast_fu_482_p1;
reg  signed [63:0] sext_ln1273_cast_reg_6613;
reg   [0:0] icmp_ln24_reg_6618;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter1_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter2_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter3_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter4_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter5_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter6_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter7_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter8_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter9_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter10_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter11_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter12_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter13_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter14_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter15_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter16_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter17_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter18_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter19_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter20_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter21_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter22_reg;
reg   [0:0] icmp_ln24_reg_6618_pp0_iter23_reg;
wire   [1:0] trunc_ln25_fu_526_p1;
reg   [1:0] trunc_ln25_reg_6622;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter1_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter2_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter3_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter4_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter5_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter6_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter7_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter8_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter9_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter10_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter11_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter12_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter13_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter14_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter15_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter16_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter17_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter18_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter19_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter20_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter21_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter22_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter23_reg;
reg   [1:0] trunc_ln25_reg_6622_pp0_iter24_reg;
wire   [31:0] tmp_3_fu_530_p6;
reg  signed [31:0] tmp_3_reg_6651;
wire   [31:0] tmp_fu_544_p6;
reg  signed [31:0] tmp_reg_6656;
wire   [63:0] mul_ln1273_fu_566_p2;
reg   [63:0] mul_ln1273_reg_6661;
reg   [0:0] tmp_73_reg_6666;
reg   [31:0] trunc_ln1_reg_6672;
reg   [0:0] tmp_74_reg_6677;
reg   [0:0] tmp_75_reg_6682;
reg   [14:0] tmp_1_reg_6687;
reg   [15:0] tmp_2_reg_6692;
wire   [63:0] mul_ln1273_1_fu_628_p2;
reg   [63:0] mul_ln1273_1_reg_6698;
reg   [0:0] tmp_80_reg_6703;
reg   [0:0] tmp_80_reg_6703_pp0_iter2_reg;
wire   [31:0] tmp_6_fu_641_p6;
reg  signed [31:0] tmp_6_reg_6708;
wire   [63:0] add_ln1347_fu_817_p2;
reg   [63:0] add_ln1347_reg_6713;
reg   [0:0] tmp_78_reg_6718;
reg   [31:0] trunc_ln818_1_reg_6724;
reg   [0:0] tmp_79_reg_6729;
reg   [14:0] tmp_4_reg_6734;
reg   [15:0] tmp_5_reg_6739;
wire   [63:0] mul_ln1273_3_fu_871_p2;
reg   [63:0] mul_ln1273_3_reg_6745;
reg   [0:0] tmp_85_reg_6750;
reg   [0:0] tmp_85_reg_6750_pp0_iter3_reg;
wire   [31:0] tmp_9_fu_884_p6;
reg  signed [31:0] tmp_9_reg_6755;
wire   [63:0] add_ln1347_1_fu_1060_p2;
reg   [63:0] add_ln1347_1_reg_6760;
reg   [0:0] tmp_83_reg_6765;
reg   [31:0] trunc_ln818_3_reg_6771;
reg   [0:0] tmp_84_reg_6776;
reg   [14:0] tmp_7_reg_6781;
reg   [15:0] tmp_8_reg_6786;
wire   [63:0] mul_ln1273_6_fu_1114_p2;
reg   [63:0] mul_ln1273_6_reg_6792;
reg   [0:0] tmp_90_reg_6797;
reg   [0:0] tmp_90_reg_6797_pp0_iter4_reg;
wire   [31:0] tmp_s_fu_1127_p6;
reg  signed [31:0] tmp_s_reg_6802;
wire   [63:0] add_ln1347_3_fu_1303_p2;
reg   [63:0] add_ln1347_3_reg_6807;
reg   [0:0] tmp_88_reg_6812;
reg   [31:0] trunc_ln818_6_reg_6818;
reg   [0:0] tmp_89_reg_6823;
reg   [14:0] tmp_10_reg_6828;
reg   [15:0] tmp_11_reg_6833;
wire   [63:0] mul_ln1273_7_fu_1357_p2;
reg   [63:0] mul_ln1273_7_reg_6839;
reg   [0:0] tmp_95_reg_6844;
reg   [0:0] tmp_95_reg_6844_pp0_iter5_reg;
wire   [31:0] tmp_14_fu_1370_p6;
reg  signed [31:0] tmp_14_reg_6849;
wire   [63:0] add_ln1347_4_fu_1546_p2;
reg   [63:0] add_ln1347_4_reg_6854;
reg   [0:0] tmp_93_reg_6859;
reg   [31:0] trunc_ln818_9_reg_6865;
reg   [0:0] tmp_94_reg_6870;
reg   [14:0] tmp_12_reg_6875;
reg   [15:0] tmp_13_reg_6880;
wire   [63:0] mul_ln1273_8_fu_1600_p2;
reg   [63:0] mul_ln1273_8_reg_6886;
reg   [0:0] tmp_100_reg_6891;
reg   [0:0] tmp_100_reg_6891_pp0_iter6_reg;
wire   [31:0] tmp_17_fu_1613_p6;
reg  signed [31:0] tmp_17_reg_6896;
wire   [63:0] add_ln1347_5_fu_1789_p2;
reg   [63:0] add_ln1347_5_reg_6901;
reg   [0:0] tmp_98_reg_6906;
reg   [31:0] trunc_ln818_s_reg_6912;
reg   [0:0] tmp_99_reg_6917;
reg   [14:0] tmp_15_reg_6922;
reg   [15:0] tmp_16_reg_6927;
wire   [63:0] mul_ln1273_9_fu_1843_p2;
reg   [63:0] mul_ln1273_9_reg_6933;
reg   [0:0] tmp_105_reg_6938;
reg   [0:0] tmp_105_reg_6938_pp0_iter7_reg;
wire   [31:0] tmp_20_fu_1856_p6;
reg  signed [31:0] tmp_20_reg_6943;
wire   [63:0] add_ln1347_6_fu_2032_p2;
reg   [63:0] add_ln1347_6_reg_6948;
reg   [0:0] tmp_103_reg_6953;
reg   [31:0] trunc_ln818_2_reg_6959;
reg   [0:0] tmp_104_reg_6964;
reg   [14:0] tmp_18_reg_6969;
reg   [15:0] tmp_19_reg_6974;
wire   [63:0] mul_ln1273_10_fu_2086_p2;
reg   [63:0] mul_ln1273_10_reg_6980;
reg   [0:0] tmp_110_reg_6985;
reg   [0:0] tmp_110_reg_6985_pp0_iter8_reg;
wire   [31:0] tmp_23_fu_2099_p6;
reg  signed [31:0] tmp_23_reg_6990;
wire   [63:0] add_ln1347_7_fu_2275_p2;
reg   [63:0] add_ln1347_7_reg_6995;
reg   [0:0] tmp_108_reg_7000;
reg   [31:0] trunc_ln818_4_reg_7006;
reg   [0:0] tmp_109_reg_7011;
reg   [14:0] tmp_21_reg_7016;
reg   [15:0] tmp_22_reg_7021;
wire   [63:0] mul_ln1273_11_fu_2329_p2;
reg   [63:0] mul_ln1273_11_reg_7027;
reg   [0:0] tmp_115_reg_7032;
reg   [0:0] tmp_115_reg_7032_pp0_iter9_reg;
wire   [31:0] tmp_26_fu_2342_p6;
reg  signed [31:0] tmp_26_reg_7037;
wire   [63:0] add_ln1347_8_fu_2518_p2;
reg   [63:0] add_ln1347_8_reg_7042;
reg   [0:0] tmp_113_reg_7047;
reg   [31:0] trunc_ln818_5_reg_7053;
reg   [0:0] tmp_114_reg_7058;
reg   [14:0] tmp_24_reg_7063;
reg   [15:0] tmp_25_reg_7068;
wire   [63:0] mul_ln1273_12_fu_2572_p2;
reg   [63:0] mul_ln1273_12_reg_7074;
reg   [0:0] tmp_120_reg_7079;
reg   [0:0] tmp_120_reg_7079_pp0_iter10_reg;
wire   [31:0] tmp_29_fu_2585_p6;
reg  signed [31:0] tmp_29_reg_7084;
wire   [63:0] add_ln1347_9_fu_2761_p2;
reg   [63:0] add_ln1347_9_reg_7089;
reg   [0:0] tmp_118_reg_7094;
reg   [31:0] trunc_ln818_7_reg_7100;
reg   [0:0] tmp_119_reg_7105;
reg   [14:0] tmp_27_reg_7110;
reg   [15:0] tmp_28_reg_7115;
wire   [63:0] mul_ln1273_13_fu_2815_p2;
reg   [63:0] mul_ln1273_13_reg_7121;
reg   [0:0] tmp_125_reg_7126;
reg   [0:0] tmp_125_reg_7126_pp0_iter11_reg;
wire   [31:0] tmp_32_fu_2828_p6;
reg  signed [31:0] tmp_32_reg_7131;
wire   [63:0] add_ln1347_10_fu_3004_p2;
reg   [63:0] add_ln1347_10_reg_7136;
reg   [0:0] tmp_123_reg_7141;
reg   [31:0] trunc_ln818_8_reg_7147;
reg   [0:0] tmp_124_reg_7152;
reg   [14:0] tmp_30_reg_7157;
reg   [15:0] tmp_31_reg_7162;
wire   [63:0] mul_ln1273_14_fu_3058_p2;
reg   [63:0] mul_ln1273_14_reg_7168;
reg   [0:0] tmp_130_reg_7173;
reg   [0:0] tmp_130_reg_7173_pp0_iter12_reg;
wire   [31:0] tmp_35_fu_3071_p6;
reg  signed [31:0] tmp_35_reg_7178;
wire   [63:0] add_ln1347_11_fu_3247_p2;
reg   [63:0] add_ln1347_11_reg_7183;
reg   [0:0] tmp_128_reg_7188;
reg   [31:0] trunc_ln818_10_reg_7194;
reg   [0:0] tmp_129_reg_7199;
reg   [14:0] tmp_33_reg_7204;
reg   [15:0] tmp_34_reg_7209;
wire   [63:0] mul_ln1273_15_fu_3301_p2;
reg   [63:0] mul_ln1273_15_reg_7215;
reg   [0:0] tmp_135_reg_7220;
reg   [0:0] tmp_135_reg_7220_pp0_iter13_reg;
wire   [31:0] tmp_38_fu_3314_p6;
reg  signed [31:0] tmp_38_reg_7225;
wire   [63:0] add_ln1347_12_fu_3490_p2;
reg   [63:0] add_ln1347_12_reg_7230;
reg   [0:0] tmp_133_reg_7235;
reg   [31:0] trunc_ln818_11_reg_7241;
reg   [0:0] tmp_134_reg_7246;
reg   [14:0] tmp_36_reg_7251;
reg   [15:0] tmp_37_reg_7256;
wire   [63:0] mul_ln1273_16_fu_3544_p2;
reg   [63:0] mul_ln1273_16_reg_7262;
reg   [0:0] tmp_140_reg_7267;
reg   [0:0] tmp_140_reg_7267_pp0_iter14_reg;
wire   [31:0] tmp_41_fu_3557_p6;
reg  signed [31:0] tmp_41_reg_7272;
wire   [63:0] add_ln1347_13_fu_3733_p2;
reg   [63:0] add_ln1347_13_reg_7277;
reg   [0:0] tmp_138_reg_7282;
reg   [31:0] trunc_ln818_12_reg_7288;
reg   [0:0] tmp_139_reg_7293;
reg   [14:0] tmp_39_reg_7298;
reg   [15:0] tmp_40_reg_7303;
wire   [63:0] mul_ln1273_17_fu_3787_p2;
reg   [63:0] mul_ln1273_17_reg_7309;
reg   [0:0] tmp_145_reg_7314;
reg   [0:0] tmp_145_reg_7314_pp0_iter15_reg;
wire   [31:0] tmp_44_fu_3800_p6;
reg  signed [31:0] tmp_44_reg_7319;
wire   [63:0] add_ln1347_14_fu_3976_p2;
reg   [63:0] add_ln1347_14_reg_7324;
reg   [0:0] tmp_143_reg_7329;
reg   [31:0] trunc_ln818_13_reg_7335;
reg   [0:0] tmp_144_reg_7340;
reg   [14:0] tmp_42_reg_7345;
reg   [15:0] tmp_43_reg_7350;
wire   [63:0] mul_ln1273_18_fu_4030_p2;
reg   [63:0] mul_ln1273_18_reg_7356;
reg   [0:0] tmp_150_reg_7361;
reg   [0:0] tmp_150_reg_7361_pp0_iter16_reg;
wire   [31:0] tmp_47_fu_4043_p6;
reg  signed [31:0] tmp_47_reg_7366;
wire   [63:0] add_ln1347_15_fu_4219_p2;
reg   [63:0] add_ln1347_15_reg_7371;
reg   [0:0] tmp_148_reg_7376;
reg   [31:0] trunc_ln818_14_reg_7382;
reg   [0:0] tmp_149_reg_7387;
reg   [14:0] tmp_45_reg_7392;
reg   [15:0] tmp_46_reg_7397;
wire   [63:0] mul_ln1273_19_fu_4273_p2;
reg   [63:0] mul_ln1273_19_reg_7403;
reg   [0:0] tmp_155_reg_7408;
reg   [0:0] tmp_155_reg_7408_pp0_iter17_reg;
wire   [31:0] tmp_50_fu_4286_p6;
reg  signed [31:0] tmp_50_reg_7413;
wire   [63:0] add_ln1347_16_fu_4462_p2;
reg   [63:0] add_ln1347_16_reg_7418;
reg   [0:0] tmp_153_reg_7423;
reg   [31:0] trunc_ln818_15_reg_7429;
reg   [0:0] tmp_154_reg_7434;
reg   [14:0] tmp_48_reg_7439;
reg   [15:0] tmp_49_reg_7444;
wire   [63:0] mul_ln1273_20_fu_4516_p2;
reg   [63:0] mul_ln1273_20_reg_7450;
reg   [0:0] tmp_160_reg_7455;
reg   [0:0] tmp_160_reg_7455_pp0_iter18_reg;
wire   [31:0] tmp_53_fu_4529_p6;
reg  signed [31:0] tmp_53_reg_7460;
wire   [63:0] add_ln1347_17_fu_4705_p2;
reg   [63:0] add_ln1347_17_reg_7465;
reg   [0:0] tmp_158_reg_7470;
reg   [31:0] trunc_ln818_16_reg_7476;
reg   [0:0] tmp_159_reg_7481;
reg   [14:0] tmp_51_reg_7486;
reg   [15:0] tmp_52_reg_7491;
wire   [63:0] mul_ln1273_21_fu_4759_p2;
reg   [63:0] mul_ln1273_21_reg_7497;
reg   [0:0] tmp_165_reg_7502;
reg   [0:0] tmp_165_reg_7502_pp0_iter19_reg;
wire   [31:0] tmp_56_fu_4772_p6;
reg  signed [31:0] tmp_56_reg_7507;
wire   [63:0] add_ln1347_18_fu_4948_p2;
reg   [63:0] add_ln1347_18_reg_7512;
reg   [0:0] tmp_163_reg_7517;
reg   [31:0] trunc_ln818_17_reg_7523;
reg   [0:0] tmp_164_reg_7528;
reg   [14:0] tmp_54_reg_7533;
reg   [15:0] tmp_55_reg_7538;
wire   [63:0] mul_ln1273_22_fu_5002_p2;
reg   [63:0] mul_ln1273_22_reg_7544;
reg   [0:0] tmp_170_reg_7549;
reg   [0:0] tmp_170_reg_7549_pp0_iter20_reg;
wire   [31:0] tmp_59_fu_5015_p6;
reg  signed [31:0] tmp_59_reg_7554;
wire   [63:0] add_ln1347_19_fu_5191_p2;
reg   [63:0] add_ln1347_19_reg_7559;
reg   [0:0] tmp_168_reg_7564;
reg   [31:0] trunc_ln818_18_reg_7570;
reg   [0:0] tmp_169_reg_7575;
reg   [14:0] tmp_57_reg_7580;
reg   [15:0] tmp_58_reg_7585;
wire   [63:0] mul_ln1273_23_fu_5245_p2;
reg   [63:0] mul_ln1273_23_reg_7591;
reg   [0:0] tmp_175_reg_7596;
reg   [0:0] tmp_175_reg_7596_pp0_iter21_reg;
wire   [31:0] tmp_62_fu_5258_p6;
reg  signed [31:0] tmp_62_reg_7601;
wire   [63:0] add_ln1347_20_fu_5434_p2;
reg   [63:0] add_ln1347_20_reg_7606;
reg   [0:0] tmp_173_reg_7611;
reg   [31:0] trunc_ln818_19_reg_7617;
reg   [0:0] tmp_174_reg_7622;
reg   [14:0] tmp_60_reg_7627;
reg   [15:0] tmp_61_reg_7632;
wire   [63:0] mul_ln1273_24_fu_5488_p2;
reg   [63:0] mul_ln1273_24_reg_7638;
reg   [0:0] tmp_180_reg_7643;
reg   [0:0] tmp_180_reg_7643_pp0_iter22_reg;
wire   [31:0] tmp_65_fu_5501_p6;
reg  signed [31:0] tmp_65_reg_7648;
wire   [63:0] add_ln1347_21_fu_5677_p2;
reg   [63:0] add_ln1347_21_reg_7653;
reg   [0:0] tmp_178_reg_7658;
reg   [31:0] trunc_ln818_20_reg_7664;
reg   [0:0] tmp_179_reg_7669;
reg   [14:0] tmp_63_reg_7674;
reg   [15:0] tmp_64_reg_7679;
wire   [63:0] mul_ln1273_25_fu_5731_p2;
reg   [63:0] mul_ln1273_25_reg_7685;
reg   [0:0] tmp_185_reg_7690;
reg   [0:0] tmp_185_reg_7690_pp0_iter23_reg;
wire   [31:0] tmp_68_fu_5744_p6;
reg  signed [31:0] tmp_68_reg_7695;
wire   [63:0] add_ln1347_22_fu_5920_p2;
reg   [63:0] add_ln1347_22_reg_7700;
reg   [0:0] tmp_183_reg_7705;
reg   [31:0] trunc_ln818_21_reg_7711;
reg   [0:0] tmp_184_reg_7716;
reg   [14:0] tmp_66_reg_7721;
reg   [15:0] tmp_67_reg_7726;
wire   [63:0] mul_ln1273_26_fu_5974_p2;
reg   [63:0] mul_ln1273_26_reg_7732;
reg   [0:0] tmp_190_reg_7737;
reg   [0:0] tmp_190_reg_7737_pp0_iter24_reg;
wire   [63:0] add_ln1347_23_fu_6150_p2;
reg   [63:0] add_ln1347_23_reg_7742;
reg   [0:0] tmp_188_reg_7747;
reg   [31:0] trunc_ln818_22_reg_7753;
reg   [0:0] tmp_189_reg_7758;
reg   [14:0] tmp_69_reg_7763;
reg   [15:0] tmp_70_reg_7768;
reg   [2:0] i_2_fu_174;
wire   [2:0] add_ln24_fu_520_p2;
wire    ap_loop_init;
reg   [2:0] ap_sig_allocacmp_i;
wire    ap_block_pp0_stage0;
reg   [31:0] temp1_V_3_2_fu_178;
wire   [31:0] temp1_V_3_8_fu_6415_p3;
reg   [31:0] temp1_V_3_3_fu_182;
wire   [31:0] temp1_V_3_7_fu_6407_p3;
reg   [31:0] temp1_V_3_4_fu_186;
wire   [31:0] temp1_V_3_6_fu_6399_p3;
reg   [31:0] temp1_V_3_1_fu_190;
wire   [31:0] temp1_V_3_fu_6391_p3;
wire    ap_block_pp0_stage0_01001;
wire  signed [31:0] mul_ln1273_fu_566_p0;
wire  signed [31:0] mul_ln1273_1_fu_628_p0;
wire   [31:0] zext_ln377_fu_654_p1;
wire   [31:0] add_ln377_fu_657_p2;
wire   [0:0] tmp_76_fu_662_p3;
wire   [0:0] xor_ln896_fu_670_p2;
wire   [0:0] and_ln378_fu_676_p2;
wire   [0:0] icmp_ln1019_1_fu_686_p2;
wire   [0:0] icmp_ln878_fu_691_p2;
wire   [0:0] tmp_77_fu_704_p3;
wire   [0:0] icmp_ln1019_fu_681_p2;
wire   [0:0] xor_ln890_fu_711_p2;
wire   [0:0] and_ln890_fu_717_p2;
wire   [0:0] select_ln888_fu_696_p3;
wire   [0:0] xor_ln895_2_fu_737_p2;
wire   [0:0] or_ln895_fu_743_p2;
wire   [0:0] xor_ln895_3_fu_749_p2;
wire   [0:0] select_ln890_fu_723_p3;
wire   [0:0] xor_ln896_1_fu_760_p2;
wire   [0:0] and_ln891_fu_731_p2;
wire   [0:0] or_ln896_fu_766_p2;
wire   [0:0] xor_ln896_20_fu_772_p2;
wire   [0:0] and_ln895_fu_754_p2;
wire   [0:0] and_ln896_fu_778_p2;
wire   [0:0] or_ln346_fu_783_p2;
wire   [31:0] select_ln346_2_fu_789_p3;
wire   [31:0] select_ln346_3_fu_797_p3;
wire   [47:0] shl_ln_fu_805_p3;
wire  signed [63:0] sext_ln813_3_fu_813_p1;
wire  signed [31:0] mul_ln1273_3_fu_871_p0;
wire   [31:0] zext_ln377_1_fu_897_p1;
wire   [31:0] add_ln377_1_fu_900_p2;
wire   [0:0] tmp_81_fu_905_p3;
wire   [0:0] xor_ln896_2_fu_913_p2;
wire   [0:0] and_ln378_1_fu_919_p2;
wire   [0:0] icmp_ln1019_3_fu_929_p2;
wire   [0:0] icmp_ln878_1_fu_934_p2;
wire   [0:0] tmp_82_fu_947_p3;
wire   [0:0] icmp_ln1019_2_fu_924_p2;
wire   [0:0] xor_ln890_7_fu_954_p2;
wire   [0:0] and_ln890_1_fu_960_p2;
wire   [0:0] select_ln888_1_fu_939_p3;
wire   [0:0] xor_ln895_4_fu_980_p2;
wire   [0:0] or_ln895_1_fu_986_p2;
wire   [0:0] xor_ln895_5_fu_992_p2;
wire   [0:0] select_ln890_1_fu_966_p3;
wire   [0:0] xor_ln896_4_fu_1003_p2;
wire   [0:0] and_ln891_1_fu_974_p2;
wire   [0:0] or_ln896_1_fu_1009_p2;
wire   [0:0] xor_ln896_23_fu_1015_p2;
wire   [0:0] and_ln895_1_fu_997_p2;
wire   [0:0] and_ln896_1_fu_1021_p2;
wire   [0:0] or_ln346_1_fu_1026_p2;
wire   [31:0] select_ln346_4_fu_1032_p3;
wire   [31:0] select_ln346_5_fu_1040_p3;
wire   [47:0] shl_ln838_1_fu_1048_p3;
wire  signed [63:0] sext_ln813_4_fu_1056_p1;
wire  signed [31:0] mul_ln1273_6_fu_1114_p0;
wire   [31:0] zext_ln377_2_fu_1140_p1;
wire   [31:0] add_ln377_3_fu_1143_p2;
wire   [0:0] tmp_86_fu_1148_p3;
wire   [0:0] xor_ln896_5_fu_1156_p2;
wire   [0:0] and_ln378_3_fu_1162_p2;
wire   [0:0] icmp_ln1019_7_fu_1172_p2;
wire   [0:0] icmp_ln878_3_fu_1177_p2;
wire   [0:0] tmp_87_fu_1190_p3;
wire   [0:0] icmp_ln1019_6_fu_1167_p2;
wire   [0:0] xor_ln890_8_fu_1197_p2;
wire   [0:0] and_ln890_2_fu_1203_p2;
wire   [0:0] select_ln888_3_fu_1182_p3;
wire   [0:0] xor_ln895_10_fu_1223_p2;
wire   [0:0] or_ln895_17_fu_1229_p2;
wire   [0:0] xor_ln895_11_fu_1235_p2;
wire   [0:0] select_ln890_3_fu_1209_p3;
wire   [0:0] xor_ln896_9_fu_1246_p2;
wire   [0:0] and_ln891_24_fu_1217_p2;
wire   [0:0] or_ln896_18_fu_1252_p2;
wire   [0:0] xor_ln896_24_fu_1258_p2;
wire   [0:0] and_ln895_3_fu_1240_p2;
wire   [0:0] and_ln896_3_fu_1264_p2;
wire   [0:0] or_ln346_3_fu_1269_p2;
wire   [31:0] select_ln346_6_fu_1275_p3;
wire   [31:0] select_ln346_7_fu_1283_p3;
wire   [47:0] shl_ln838_3_fu_1291_p3;
wire  signed [63:0] sext_ln813_5_fu_1299_p1;
wire  signed [31:0] mul_ln1273_7_fu_1357_p0;
wire   [31:0] zext_ln377_3_fu_1383_p1;
wire   [31:0] add_ln377_6_fu_1386_p2;
wire   [0:0] tmp_91_fu_1391_p3;
wire   [0:0] xor_ln896_10_fu_1399_p2;
wire   [0:0] and_ln378_6_fu_1405_p2;
wire   [0:0] icmp_ln1019_9_fu_1415_p2;
wire   [0:0] icmp_ln878_4_fu_1420_p2;
wire   [0:0] tmp_92_fu_1433_p3;
wire   [0:0] icmp_ln1019_8_fu_1410_p2;
wire   [0:0] xor_ln890_9_fu_1440_p2;
wire   [0:0] and_ln890_3_fu_1446_p2;
wire   [0:0] select_ln888_4_fu_1425_p3;
wire   [0:0] xor_ln895_fu_1466_p2;
wire   [0:0] or_ln895_3_fu_1472_p2;
wire   [0:0] xor_ln895_14_fu_1478_p2;
wire   [0:0] select_ln890_4_fu_1452_p3;
wire   [0:0] xor_ln896_15_fu_1489_p2;
wire   [0:0] and_ln891_3_fu_1460_p2;
wire   [0:0] or_ln896_3_fu_1495_p2;
wire   [0:0] xor_ln896_25_fu_1501_p2;
wire   [0:0] and_ln895_6_fu_1483_p2;
wire   [0:0] and_ln896_6_fu_1507_p2;
wire   [0:0] or_ln346_6_fu_1512_p2;
wire   [31:0] select_ln346_8_fu_1518_p3;
wire   [31:0] select_ln346_9_fu_1526_p3;
wire   [47:0] shl_ln838_6_fu_1534_p3;
wire  signed [63:0] sext_ln813_6_fu_1542_p1;
wire  signed [31:0] mul_ln1273_8_fu_1600_p0;
wire   [31:0] zext_ln377_4_fu_1626_p1;
wire   [31:0] add_ln377_7_fu_1629_p2;
wire   [0:0] tmp_96_fu_1634_p3;
wire   [0:0] xor_ln896_16_fu_1642_p2;
wire   [0:0] and_ln378_7_fu_1648_p2;
wire   [0:0] icmp_ln1019_11_fu_1658_p2;
wire   [0:0] icmp_ln878_5_fu_1663_p2;
wire   [0:0] tmp_97_fu_1676_p3;
wire   [0:0] icmp_ln1019_10_fu_1653_p2;
wire   [0:0] xor_ln890_10_fu_1683_p2;
wire   [0:0] and_ln890_4_fu_1689_p2;
wire   [0:0] select_ln888_5_fu_1668_p3;
wire   [0:0] xor_ln895_15_fu_1709_p2;
wire   [0:0] or_ln895_4_fu_1715_p2;
wire   [0:0] xor_ln895_16_fu_1721_p2;
wire   [0:0] select_ln890_5_fu_1695_p3;
wire   [0:0] xor_ln896_21_fu_1732_p2;
wire   [0:0] and_ln891_4_fu_1703_p2;
wire   [0:0] or_ln896_4_fu_1738_p2;
wire   [0:0] xor_ln896_28_fu_1744_p2;
wire   [0:0] and_ln895_7_fu_1726_p2;
wire   [0:0] and_ln896_7_fu_1750_p2;
wire   [0:0] or_ln346_7_fu_1755_p2;
wire   [31:0] select_ln346_10_fu_1761_p3;
wire   [31:0] select_ln346_11_fu_1769_p3;
wire   [47:0] shl_ln838_9_fu_1777_p3;
wire  signed [63:0] sext_ln813_7_fu_1785_p1;
wire  signed [31:0] mul_ln1273_9_fu_1843_p0;
wire   [31:0] zext_ln377_5_fu_1869_p1;
wire   [31:0] add_ln377_8_fu_1872_p2;
wire   [0:0] tmp_101_fu_1877_p3;
wire   [0:0] xor_ln896_22_fu_1885_p2;
wire   [0:0] and_ln378_8_fu_1891_p2;
wire   [0:0] icmp_ln1019_13_fu_1901_p2;
wire   [0:0] icmp_ln878_6_fu_1906_p2;
wire   [0:0] tmp_102_fu_1919_p3;
wire   [0:0] icmp_ln1019_12_fu_1896_p2;
wire   [0:0] xor_ln890_11_fu_1926_p2;
wire   [0:0] and_ln890_5_fu_1932_p2;
wire   [0:0] select_ln888_6_fu_1911_p3;
wire   [0:0] xor_ln895_17_fu_1952_p2;
wire   [0:0] or_ln895_5_fu_1958_p2;
wire   [0:0] xor_ln895_18_fu_1964_p2;
wire   [0:0] select_ln890_6_fu_1938_p3;
wire   [0:0] xor_ln896_26_fu_1975_p2;
wire   [0:0] and_ln891_5_fu_1946_p2;
wire   [0:0] or_ln896_5_fu_1981_p2;
wire   [0:0] xor_ln896_64_fu_1987_p2;
wire   [0:0] and_ln895_8_fu_1969_p2;
wire   [0:0] and_ln896_8_fu_1993_p2;
wire   [0:0] or_ln346_8_fu_1998_p2;
wire   [31:0] select_ln346_12_fu_2004_p3;
wire   [31:0] select_ln346_13_fu_2012_p3;
wire   [47:0] shl_ln838_s_fu_2020_p3;
wire  signed [63:0] sext_ln813_8_fu_2028_p1;
wire  signed [31:0] mul_ln1273_10_fu_2086_p0;
wire   [31:0] zext_ln377_6_fu_2112_p1;
wire   [31:0] add_ln377_9_fu_2115_p2;
wire   [0:0] tmp_106_fu_2120_p3;
wire   [0:0] xor_ln896_27_fu_2128_p2;
wire   [0:0] and_ln378_9_fu_2134_p2;
wire   [0:0] icmp_ln1019_15_fu_2144_p2;
wire   [0:0] icmp_ln878_7_fu_2149_p2;
wire   [0:0] tmp_107_fu_2162_p3;
wire   [0:0] icmp_ln1019_14_fu_2139_p2;
wire   [0:0] xor_ln890_12_fu_2169_p2;
wire   [0:0] and_ln890_6_fu_2175_p2;
wire   [0:0] select_ln888_7_fu_2154_p3;
wire   [0:0] xor_ln895_19_fu_2195_p2;
wire   [0:0] or_ln895_6_fu_2201_p2;
wire   [0:0] xor_ln895_20_fu_2207_p2;
wire   [0:0] select_ln890_7_fu_2181_p3;
wire   [0:0] xor_ln896_29_fu_2218_p2;
wire   [0:0] and_ln891_6_fu_2189_p2;
wire   [0:0] or_ln896_6_fu_2224_p2;
wire   [0:0] xor_ln896_65_fu_2230_p2;
wire   [0:0] and_ln895_9_fu_2212_p2;
wire   [0:0] and_ln896_9_fu_2236_p2;
wire   [0:0] or_ln346_9_fu_2241_p2;
wire   [31:0] select_ln346_14_fu_2247_p3;
wire   [31:0] select_ln346_fu_2255_p3;
wire   [47:0] shl_ln838_2_fu_2263_p3;
wire  signed [63:0] sext_ln813_fu_2271_p1;
wire  signed [31:0] mul_ln1273_11_fu_2329_p0;
wire   [31:0] zext_ln377_7_fu_2355_p1;
wire   [31:0] add_ln377_10_fu_2358_p2;
wire   [0:0] tmp_111_fu_2363_p3;
wire   [0:0] xor_ln896_30_fu_2371_p2;
wire   [0:0] and_ln378_10_fu_2377_p2;
wire   [0:0] icmp_ln1019_17_fu_2387_p2;
wire   [0:0] icmp_ln878_8_fu_2392_p2;
wire   [0:0] tmp_112_fu_2405_p3;
wire   [0:0] icmp_ln1019_16_fu_2382_p2;
wire   [0:0] xor_ln890_13_fu_2412_p2;
wire   [0:0] and_ln890_7_fu_2418_p2;
wire   [0:0] select_ln888_8_fu_2397_p3;
wire   [0:0] xor_ln895_21_fu_2438_p2;
wire   [0:0] or_ln895_7_fu_2444_p2;
wire   [0:0] xor_ln895_22_fu_2450_p2;
wire   [0:0] select_ln890_8_fu_2424_p3;
wire   [0:0] xor_ln896_31_fu_2461_p2;
wire   [0:0] and_ln891_7_fu_2432_p2;
wire   [0:0] or_ln896_7_fu_2467_p2;
wire   [0:0] xor_ln896_66_fu_2473_p2;
wire   [0:0] and_ln895_10_fu_2455_p2;
wire   [0:0] and_ln896_10_fu_2479_p2;
wire   [0:0] or_ln346_10_fu_2484_p2;
wire   [31:0] select_ln346_15_fu_2490_p3;
wire   [31:0] select_ln346_16_fu_2498_p3;
wire   [47:0] shl_ln838_4_fu_2506_p3;
wire  signed [63:0] sext_ln813_9_fu_2514_p1;
wire  signed [31:0] mul_ln1273_12_fu_2572_p0;
wire   [31:0] zext_ln377_8_fu_2598_p1;
wire   [31:0] add_ln377_11_fu_2601_p2;
wire   [0:0] tmp_116_fu_2606_p3;
wire   [0:0] xor_ln896_32_fu_2614_p2;
wire   [0:0] and_ln378_11_fu_2620_p2;
wire   [0:0] icmp_ln1019_19_fu_2630_p2;
wire   [0:0] icmp_ln878_9_fu_2635_p2;
wire   [0:0] tmp_117_fu_2648_p3;
wire   [0:0] icmp_ln1019_18_fu_2625_p2;
wire   [0:0] xor_ln890_14_fu_2655_p2;
wire   [0:0] and_ln890_8_fu_2661_p2;
wire   [0:0] select_ln888_9_fu_2640_p3;
wire   [0:0] xor_ln895_23_fu_2681_p2;
wire   [0:0] or_ln895_8_fu_2687_p2;
wire   [0:0] xor_ln895_24_fu_2693_p2;
wire   [0:0] select_ln890_9_fu_2667_p3;
wire   [0:0] xor_ln896_33_fu_2704_p2;
wire   [0:0] and_ln891_8_fu_2675_p2;
wire   [0:0] or_ln896_8_fu_2710_p2;
wire   [0:0] xor_ln896_67_fu_2716_p2;
wire   [0:0] and_ln895_11_fu_2698_p2;
wire   [0:0] and_ln896_11_fu_2722_p2;
wire   [0:0] or_ln346_11_fu_2727_p2;
wire   [31:0] select_ln346_17_fu_2733_p3;
wire   [31:0] select_ln346_18_fu_2741_p3;
wire   [47:0] shl_ln838_5_fu_2749_p3;
wire  signed [63:0] sext_ln813_10_fu_2757_p1;
wire  signed [31:0] mul_ln1273_13_fu_2815_p0;
wire   [31:0] zext_ln377_9_fu_2841_p1;
wire   [31:0] add_ln377_12_fu_2844_p2;
wire   [0:0] tmp_121_fu_2849_p3;
wire   [0:0] xor_ln896_34_fu_2857_p2;
wire   [0:0] and_ln378_12_fu_2863_p2;
wire   [0:0] icmp_ln1019_21_fu_2873_p2;
wire   [0:0] icmp_ln878_10_fu_2878_p2;
wire   [0:0] tmp_122_fu_2891_p3;
wire   [0:0] icmp_ln1019_20_fu_2868_p2;
wire   [0:0] xor_ln890_15_fu_2898_p2;
wire   [0:0] and_ln890_9_fu_2904_p2;
wire   [0:0] select_ln888_10_fu_2883_p3;
wire   [0:0] xor_ln895_25_fu_2924_p2;
wire   [0:0] or_ln895_9_fu_2930_p2;
wire   [0:0] xor_ln895_26_fu_2936_p2;
wire   [0:0] select_ln890_10_fu_2910_p3;
wire   [0:0] xor_ln896_35_fu_2947_p2;
wire   [0:0] and_ln891_9_fu_2918_p2;
wire   [0:0] or_ln896_9_fu_2953_p2;
wire   [0:0] xor_ln896_68_fu_2959_p2;
wire   [0:0] and_ln895_12_fu_2941_p2;
wire   [0:0] and_ln896_12_fu_2965_p2;
wire   [0:0] or_ln346_12_fu_2970_p2;
wire   [31:0] select_ln346_19_fu_2976_p3;
wire   [31:0] select_ln346_20_fu_2984_p3;
wire   [47:0] shl_ln838_7_fu_2992_p3;
wire  signed [63:0] sext_ln813_11_fu_3000_p1;
wire  signed [31:0] mul_ln1273_14_fu_3058_p0;
wire   [31:0] zext_ln377_10_fu_3084_p1;
wire   [31:0] add_ln377_13_fu_3087_p2;
wire   [0:0] tmp_126_fu_3092_p3;
wire   [0:0] xor_ln896_36_fu_3100_p2;
wire   [0:0] and_ln378_13_fu_3106_p2;
wire   [0:0] icmp_ln1019_23_fu_3116_p2;
wire   [0:0] icmp_ln878_11_fu_3121_p2;
wire   [0:0] tmp_127_fu_3134_p3;
wire   [0:0] icmp_ln1019_22_fu_3111_p2;
wire   [0:0] xor_ln890_16_fu_3141_p2;
wire   [0:0] and_ln890_10_fu_3147_p2;
wire   [0:0] select_ln888_11_fu_3126_p3;
wire   [0:0] xor_ln895_27_fu_3167_p2;
wire   [0:0] or_ln895_10_fu_3173_p2;
wire   [0:0] xor_ln895_28_fu_3179_p2;
wire   [0:0] select_ln890_11_fu_3153_p3;
wire   [0:0] xor_ln896_37_fu_3190_p2;
wire   [0:0] and_ln891_10_fu_3161_p2;
wire   [0:0] or_ln896_10_fu_3196_p2;
wire   [0:0] xor_ln896_69_fu_3202_p2;
wire   [0:0] and_ln895_13_fu_3184_p2;
wire   [0:0] and_ln896_13_fu_3208_p2;
wire   [0:0] or_ln346_13_fu_3213_p2;
wire   [31:0] select_ln346_21_fu_3219_p3;
wire   [31:0] select_ln346_22_fu_3227_p3;
wire   [47:0] shl_ln838_8_fu_3235_p3;
wire  signed [63:0] sext_ln813_12_fu_3243_p1;
wire  signed [31:0] mul_ln1273_15_fu_3301_p0;
wire   [31:0] zext_ln377_11_fu_3327_p1;
wire   [31:0] add_ln377_14_fu_3330_p2;
wire   [0:0] tmp_131_fu_3335_p3;
wire   [0:0] xor_ln896_38_fu_3343_p2;
wire   [0:0] and_ln378_14_fu_3349_p2;
wire   [0:0] icmp_ln1019_25_fu_3359_p2;
wire   [0:0] icmp_ln878_12_fu_3364_p2;
wire   [0:0] tmp_132_fu_3377_p3;
wire   [0:0] icmp_ln1019_24_fu_3354_p2;
wire   [0:0] xor_ln890_17_fu_3384_p2;
wire   [0:0] and_ln890_11_fu_3390_p2;
wire   [0:0] select_ln888_12_fu_3369_p3;
wire   [0:0] xor_ln895_29_fu_3410_p2;
wire   [0:0] or_ln895_11_fu_3416_p2;
wire   [0:0] xor_ln895_30_fu_3422_p2;
wire   [0:0] select_ln890_12_fu_3396_p3;
wire   [0:0] xor_ln896_39_fu_3433_p2;
wire   [0:0] and_ln891_11_fu_3404_p2;
wire   [0:0] or_ln896_11_fu_3439_p2;
wire   [0:0] xor_ln896_70_fu_3445_p2;
wire   [0:0] and_ln895_14_fu_3427_p2;
wire   [0:0] and_ln896_14_fu_3451_p2;
wire   [0:0] or_ln346_14_fu_3456_p2;
wire   [31:0] select_ln346_23_fu_3462_p3;
wire   [31:0] select_ln346_24_fu_3470_p3;
wire   [47:0] shl_ln838_10_fu_3478_p3;
wire  signed [63:0] sext_ln813_13_fu_3486_p1;
wire  signed [31:0] mul_ln1273_16_fu_3544_p0;
wire   [31:0] zext_ln377_12_fu_3570_p1;
wire   [31:0] add_ln377_15_fu_3573_p2;
wire   [0:0] tmp_136_fu_3578_p3;
wire   [0:0] xor_ln896_40_fu_3586_p2;
wire   [0:0] and_ln378_15_fu_3592_p2;
wire   [0:0] icmp_ln1019_27_fu_3602_p2;
wire   [0:0] icmp_ln878_13_fu_3607_p2;
wire   [0:0] tmp_137_fu_3620_p3;
wire   [0:0] icmp_ln1019_26_fu_3597_p2;
wire   [0:0] xor_ln890_18_fu_3627_p2;
wire   [0:0] and_ln890_12_fu_3633_p2;
wire   [0:0] select_ln888_13_fu_3612_p3;
wire   [0:0] xor_ln895_31_fu_3653_p2;
wire   [0:0] or_ln895_12_fu_3659_p2;
wire   [0:0] xor_ln895_32_fu_3665_p2;
wire   [0:0] select_ln890_13_fu_3639_p3;
wire   [0:0] xor_ln896_41_fu_3676_p2;
wire   [0:0] and_ln891_12_fu_3647_p2;
wire   [0:0] or_ln896_12_fu_3682_p2;
wire   [0:0] xor_ln896_71_fu_3688_p2;
wire   [0:0] and_ln895_15_fu_3670_p2;
wire   [0:0] and_ln896_15_fu_3694_p2;
wire   [0:0] or_ln346_15_fu_3699_p2;
wire   [31:0] select_ln346_25_fu_3705_p3;
wire   [31:0] select_ln346_26_fu_3713_p3;
wire   [47:0] shl_ln838_11_fu_3721_p3;
wire  signed [63:0] sext_ln813_14_fu_3729_p1;
wire  signed [31:0] mul_ln1273_17_fu_3787_p0;
wire   [31:0] zext_ln377_13_fu_3813_p1;
wire   [31:0] add_ln377_16_fu_3816_p2;
wire   [0:0] tmp_141_fu_3821_p3;
wire   [0:0] xor_ln896_42_fu_3829_p2;
wire   [0:0] and_ln378_16_fu_3835_p2;
wire   [0:0] icmp_ln1019_29_fu_3845_p2;
wire   [0:0] icmp_ln878_14_fu_3850_p2;
wire   [0:0] tmp_142_fu_3863_p3;
wire   [0:0] icmp_ln1019_28_fu_3840_p2;
wire   [0:0] xor_ln890_19_fu_3870_p2;
wire   [0:0] and_ln890_13_fu_3876_p2;
wire   [0:0] select_ln888_14_fu_3855_p3;
wire   [0:0] xor_ln895_33_fu_3896_p2;
wire   [0:0] or_ln895_13_fu_3902_p2;
wire   [0:0] xor_ln895_34_fu_3908_p2;
wire   [0:0] select_ln890_14_fu_3882_p3;
wire   [0:0] xor_ln896_43_fu_3919_p2;
wire   [0:0] and_ln891_13_fu_3890_p2;
wire   [0:0] or_ln896_13_fu_3925_p2;
wire   [0:0] xor_ln896_72_fu_3931_p2;
wire   [0:0] and_ln895_16_fu_3913_p2;
wire   [0:0] and_ln896_16_fu_3937_p2;
wire   [0:0] or_ln346_16_fu_3942_p2;
wire   [31:0] select_ln346_27_fu_3948_p3;
wire   [31:0] select_ln346_28_fu_3956_p3;
wire   [47:0] shl_ln838_12_fu_3964_p3;
wire  signed [63:0] sext_ln813_15_fu_3972_p1;
wire  signed [31:0] mul_ln1273_18_fu_4030_p0;
wire   [31:0] zext_ln377_14_fu_4056_p1;
wire   [31:0] add_ln377_17_fu_4059_p2;
wire   [0:0] tmp_146_fu_4064_p3;
wire   [0:0] xor_ln896_44_fu_4072_p2;
wire   [0:0] and_ln378_17_fu_4078_p2;
wire   [0:0] icmp_ln1019_31_fu_4088_p2;
wire   [0:0] icmp_ln878_15_fu_4093_p2;
wire   [0:0] tmp_147_fu_4106_p3;
wire   [0:0] icmp_ln1019_30_fu_4083_p2;
wire   [0:0] xor_ln890_20_fu_4113_p2;
wire   [0:0] and_ln890_14_fu_4119_p2;
wire   [0:0] select_ln888_15_fu_4098_p3;
wire   [0:0] xor_ln895_35_fu_4139_p2;
wire   [0:0] or_ln895_14_fu_4145_p2;
wire   [0:0] xor_ln895_36_fu_4151_p2;
wire   [0:0] select_ln890_15_fu_4125_p3;
wire   [0:0] xor_ln896_45_fu_4162_p2;
wire   [0:0] and_ln891_14_fu_4133_p2;
wire   [0:0] or_ln896_14_fu_4168_p2;
wire   [0:0] xor_ln896_73_fu_4174_p2;
wire   [0:0] and_ln895_17_fu_4156_p2;
wire   [0:0] and_ln896_17_fu_4180_p2;
wire   [0:0] or_ln346_17_fu_4185_p2;
wire   [31:0] select_ln346_29_fu_4191_p3;
wire   [31:0] select_ln346_30_fu_4199_p3;
wire   [47:0] shl_ln838_13_fu_4207_p3;
wire  signed [63:0] sext_ln813_16_fu_4215_p1;
wire  signed [31:0] mul_ln1273_19_fu_4273_p0;
wire   [31:0] zext_ln377_15_fu_4299_p1;
wire   [31:0] add_ln377_18_fu_4302_p2;
wire   [0:0] tmp_151_fu_4307_p3;
wire   [0:0] xor_ln896_46_fu_4315_p2;
wire   [0:0] and_ln378_18_fu_4321_p2;
wire   [0:0] icmp_ln1019_33_fu_4331_p2;
wire   [0:0] icmp_ln878_16_fu_4336_p2;
wire   [0:0] tmp_152_fu_4349_p3;
wire   [0:0] icmp_ln1019_32_fu_4326_p2;
wire   [0:0] xor_ln890_21_fu_4356_p2;
wire   [0:0] and_ln890_15_fu_4362_p2;
wire   [0:0] select_ln888_16_fu_4341_p3;
wire   [0:0] xor_ln895_37_fu_4382_p2;
wire   [0:0] or_ln895_15_fu_4388_p2;
wire   [0:0] xor_ln895_38_fu_4394_p2;
wire   [0:0] select_ln890_16_fu_4368_p3;
wire   [0:0] xor_ln896_47_fu_4405_p2;
wire   [0:0] and_ln891_15_fu_4376_p2;
wire   [0:0] or_ln896_15_fu_4411_p2;
wire   [0:0] xor_ln896_74_fu_4417_p2;
wire   [0:0] and_ln895_18_fu_4399_p2;
wire   [0:0] and_ln896_18_fu_4423_p2;
wire   [0:0] or_ln346_18_fu_4428_p2;
wire   [31:0] select_ln346_31_fu_4434_p3;
wire   [31:0] select_ln346_32_fu_4442_p3;
wire   [47:0] shl_ln838_14_fu_4450_p3;
wire  signed [63:0] sext_ln813_17_fu_4458_p1;
wire  signed [31:0] mul_ln1273_20_fu_4516_p0;
wire   [31:0] zext_ln377_16_fu_4542_p1;
wire   [31:0] add_ln377_19_fu_4545_p2;
wire   [0:0] tmp_156_fu_4550_p3;
wire   [0:0] xor_ln896_48_fu_4558_p2;
wire   [0:0] and_ln378_19_fu_4564_p2;
wire   [0:0] icmp_ln1019_35_fu_4574_p2;
wire   [0:0] icmp_ln878_17_fu_4579_p2;
wire   [0:0] tmp_157_fu_4592_p3;
wire   [0:0] icmp_ln1019_34_fu_4569_p2;
wire   [0:0] xor_ln890_22_fu_4599_p2;
wire   [0:0] and_ln890_16_fu_4605_p2;
wire   [0:0] select_ln888_17_fu_4584_p3;
wire   [0:0] xor_ln895_39_fu_4625_p2;
wire   [0:0] or_ln895_16_fu_4631_p2;
wire   [0:0] xor_ln895_40_fu_4637_p2;
wire   [0:0] select_ln890_17_fu_4611_p3;
wire   [0:0] xor_ln896_49_fu_4648_p2;
wire   [0:0] and_ln891_16_fu_4619_p2;
wire   [0:0] or_ln896_16_fu_4654_p2;
wire   [0:0] xor_ln896_75_fu_4660_p2;
wire   [0:0] and_ln895_19_fu_4642_p2;
wire   [0:0] and_ln896_19_fu_4666_p2;
wire   [0:0] or_ln346_19_fu_4671_p2;
wire   [31:0] select_ln346_33_fu_4677_p3;
wire   [31:0] select_ln346_34_fu_4685_p3;
wire   [47:0] shl_ln838_15_fu_4693_p3;
wire  signed [63:0] sext_ln813_18_fu_4701_p1;
wire  signed [31:0] mul_ln1273_21_fu_4759_p0;
wire   [31:0] zext_ln377_17_fu_4785_p1;
wire   [31:0] add_ln377_20_fu_4788_p2;
wire   [0:0] tmp_161_fu_4793_p3;
wire   [0:0] xor_ln896_50_fu_4801_p2;
wire   [0:0] and_ln378_20_fu_4807_p2;
wire   [0:0] icmp_ln1019_37_fu_4817_p2;
wire   [0:0] icmp_ln878_18_fu_4822_p2;
wire   [0:0] tmp_162_fu_4835_p3;
wire   [0:0] icmp_ln1019_36_fu_4812_p2;
wire   [0:0] xor_ln890_23_fu_4842_p2;
wire   [0:0] and_ln890_17_fu_4848_p2;
wire   [0:0] select_ln888_18_fu_4827_p3;
wire   [0:0] xor_ln895_41_fu_4868_p2;
wire   [0:0] or_ln895_24_fu_4874_p2;
wire   [0:0] xor_ln895_42_fu_4880_p2;
wire   [0:0] select_ln890_18_fu_4854_p3;
wire   [0:0] xor_ln896_51_fu_4891_p2;
wire   [0:0] and_ln891_17_fu_4862_p2;
wire   [0:0] or_ln896_17_fu_4897_p2;
wire   [0:0] xor_ln896_76_fu_4903_p2;
wire   [0:0] and_ln895_20_fu_4885_p2;
wire   [0:0] and_ln896_20_fu_4909_p2;
wire   [0:0] or_ln346_20_fu_4914_p2;
wire   [31:0] select_ln346_35_fu_4920_p3;
wire   [31:0] select_ln346_36_fu_4928_p3;
wire   [47:0] shl_ln838_16_fu_4936_p3;
wire  signed [63:0] sext_ln813_19_fu_4944_p1;
wire  signed [31:0] mul_ln1273_22_fu_5002_p0;
wire   [31:0] zext_ln377_18_fu_5028_p1;
wire   [31:0] add_ln377_21_fu_5031_p2;
wire   [0:0] tmp_166_fu_5036_p3;
wire   [0:0] xor_ln896_52_fu_5044_p2;
wire   [0:0] and_ln378_21_fu_5050_p2;
wire   [0:0] icmp_ln1019_39_fu_5060_p2;
wire   [0:0] icmp_ln878_19_fu_5065_p2;
wire   [0:0] tmp_167_fu_5078_p3;
wire   [0:0] icmp_ln1019_38_fu_5055_p2;
wire   [0:0] xor_ln890_24_fu_5085_p2;
wire   [0:0] and_ln890_18_fu_5091_p2;
wire   [0:0] select_ln888_19_fu_5070_p3;
wire   [0:0] xor_ln895_43_fu_5111_p2;
wire   [0:0] or_ln895_18_fu_5117_p2;
wire   [0:0] xor_ln895_44_fu_5123_p2;
wire   [0:0] select_ln890_19_fu_5097_p3;
wire   [0:0] xor_ln896_53_fu_5134_p2;
wire   [0:0] and_ln891_18_fu_5105_p2;
wire   [0:0] or_ln896_24_fu_5140_p2;
wire   [0:0] xor_ln896_77_fu_5146_p2;
wire   [0:0] and_ln895_21_fu_5128_p2;
wire   [0:0] and_ln896_21_fu_5152_p2;
wire   [0:0] or_ln346_21_fu_5157_p2;
wire   [31:0] select_ln346_37_fu_5163_p3;
wire   [31:0] select_ln346_38_fu_5171_p3;
wire   [47:0] shl_ln838_17_fu_5179_p3;
wire  signed [63:0] sext_ln813_20_fu_5187_p1;
wire  signed [31:0] mul_ln1273_23_fu_5245_p0;
wire   [31:0] zext_ln377_19_fu_5271_p1;
wire   [31:0] add_ln377_22_fu_5274_p2;
wire   [0:0] tmp_171_fu_5279_p3;
wire   [0:0] xor_ln896_54_fu_5287_p2;
wire   [0:0] and_ln378_22_fu_5293_p2;
wire   [0:0] icmp_ln1019_41_fu_5303_p2;
wire   [0:0] icmp_ln878_20_fu_5308_p2;
wire   [0:0] tmp_172_fu_5321_p3;
wire   [0:0] icmp_ln1019_40_fu_5298_p2;
wire   [0:0] xor_ln890_25_fu_5328_p2;
wire   [0:0] and_ln890_19_fu_5334_p2;
wire   [0:0] select_ln888_20_fu_5313_p3;
wire   [0:0] xor_ln895_45_fu_5354_p2;
wire   [0:0] or_ln895_19_fu_5360_p2;
wire   [0:0] xor_ln895_46_fu_5366_p2;
wire   [0:0] select_ln890_20_fu_5340_p3;
wire   [0:0] xor_ln896_55_fu_5377_p2;
wire   [0:0] and_ln891_19_fu_5348_p2;
wire   [0:0] or_ln896_19_fu_5383_p2;
wire   [0:0] xor_ln896_78_fu_5389_p2;
wire   [0:0] and_ln895_22_fu_5371_p2;
wire   [0:0] and_ln896_22_fu_5395_p2;
wire   [0:0] or_ln346_22_fu_5400_p2;
wire   [31:0] select_ln346_39_fu_5406_p3;
wire   [31:0] select_ln346_40_fu_5414_p3;
wire   [47:0] shl_ln838_18_fu_5422_p3;
wire  signed [63:0] sext_ln813_21_fu_5430_p1;
wire  signed [31:0] mul_ln1273_24_fu_5488_p0;
wire   [31:0] zext_ln377_20_fu_5514_p1;
wire   [31:0] add_ln377_23_fu_5517_p2;
wire   [0:0] tmp_176_fu_5522_p3;
wire   [0:0] xor_ln896_56_fu_5530_p2;
wire   [0:0] and_ln378_23_fu_5536_p2;
wire   [0:0] icmp_ln1019_43_fu_5546_p2;
wire   [0:0] icmp_ln878_21_fu_5551_p2;
wire   [0:0] tmp_177_fu_5564_p3;
wire   [0:0] icmp_ln1019_42_fu_5541_p2;
wire   [0:0] xor_ln890_26_fu_5571_p2;
wire   [0:0] and_ln890_20_fu_5577_p2;
wire   [0:0] select_ln888_21_fu_5556_p3;
wire   [0:0] xor_ln895_47_fu_5597_p2;
wire   [0:0] or_ln895_20_fu_5603_p2;
wire   [0:0] xor_ln895_48_fu_5609_p2;
wire   [0:0] select_ln890_21_fu_5583_p3;
wire   [0:0] xor_ln896_57_fu_5620_p2;
wire   [0:0] and_ln891_20_fu_5591_p2;
wire   [0:0] or_ln896_20_fu_5626_p2;
wire   [0:0] xor_ln896_79_fu_5632_p2;
wire   [0:0] and_ln895_23_fu_5614_p2;
wire   [0:0] and_ln896_23_fu_5638_p2;
wire   [0:0] or_ln346_23_fu_5643_p2;
wire   [31:0] select_ln346_41_fu_5649_p3;
wire   [31:0] select_ln346_42_fu_5657_p3;
wire   [47:0] shl_ln838_19_fu_5665_p3;
wire  signed [63:0] sext_ln813_22_fu_5673_p1;
wire  signed [31:0] mul_ln1273_25_fu_5731_p0;
wire   [31:0] zext_ln377_21_fu_5757_p1;
wire   [31:0] add_ln377_24_fu_5760_p2;
wire   [0:0] tmp_181_fu_5765_p3;
wire   [0:0] xor_ln896_58_fu_5773_p2;
wire   [0:0] and_ln378_24_fu_5779_p2;
wire   [0:0] icmp_ln1019_45_fu_5789_p2;
wire   [0:0] icmp_ln878_22_fu_5794_p2;
wire   [0:0] tmp_182_fu_5807_p3;
wire   [0:0] icmp_ln1019_44_fu_5784_p2;
wire   [0:0] xor_ln890_27_fu_5814_p2;
wire   [0:0] and_ln890_21_fu_5820_p2;
wire   [0:0] select_ln888_22_fu_5799_p3;
wire   [0:0] xor_ln895_49_fu_5840_p2;
wire   [0:0] or_ln895_21_fu_5846_p2;
wire   [0:0] xor_ln895_50_fu_5852_p2;
wire   [0:0] select_ln890_22_fu_5826_p3;
wire   [0:0] xor_ln896_59_fu_5863_p2;
wire   [0:0] and_ln891_21_fu_5834_p2;
wire   [0:0] or_ln896_21_fu_5869_p2;
wire   [0:0] xor_ln896_80_fu_5875_p2;
wire   [0:0] and_ln895_24_fu_5857_p2;
wire   [0:0] and_ln896_24_fu_5881_p2;
wire   [0:0] or_ln346_24_fu_5886_p2;
wire   [31:0] select_ln346_43_fu_5892_p3;
wire   [31:0] select_ln346_44_fu_5900_p3;
wire   [47:0] shl_ln838_20_fu_5908_p3;
wire  signed [63:0] sext_ln813_23_fu_5916_p1;
wire  signed [31:0] mul_ln1273_26_fu_5974_p0;
wire   [31:0] zext_ln377_22_fu_5987_p1;
wire   [31:0] add_ln377_25_fu_5990_p2;
wire   [0:0] tmp_186_fu_5995_p3;
wire   [0:0] xor_ln896_60_fu_6003_p2;
wire   [0:0] and_ln378_25_fu_6009_p2;
wire   [0:0] icmp_ln1019_47_fu_6019_p2;
wire   [0:0] icmp_ln878_23_fu_6024_p2;
wire   [0:0] tmp_187_fu_6037_p3;
wire   [0:0] icmp_ln1019_46_fu_6014_p2;
wire   [0:0] xor_ln890_28_fu_6044_p2;
wire   [0:0] and_ln890_22_fu_6050_p2;
wire   [0:0] select_ln888_23_fu_6029_p3;
wire   [0:0] xor_ln895_51_fu_6070_p2;
wire   [0:0] or_ln895_22_fu_6076_p2;
wire   [0:0] xor_ln895_52_fu_6082_p2;
wire   [0:0] select_ln890_23_fu_6056_p3;
wire   [0:0] xor_ln896_61_fu_6093_p2;
wire   [0:0] and_ln891_22_fu_6064_p2;
wire   [0:0] or_ln896_22_fu_6099_p2;
wire   [0:0] xor_ln896_81_fu_6105_p2;
wire   [0:0] and_ln895_25_fu_6087_p2;
wire   [0:0] and_ln896_25_fu_6111_p2;
wire   [0:0] or_ln346_25_fu_6116_p2;
wire   [31:0] select_ln346_45_fu_6122_p3;
wire   [31:0] select_ln346_46_fu_6130_p3;
wire   [47:0] shl_ln838_21_fu_6138_p3;
wire  signed [63:0] sext_ln813_24_fu_6146_p1;
wire   [31:0] zext_ln377_23_fu_6213_p1;
wire   [31:0] add_ln377_26_fu_6216_p2;
wire   [0:0] tmp_191_fu_6221_p3;
wire   [0:0] xor_ln896_62_fu_6229_p2;
wire   [0:0] and_ln378_26_fu_6235_p2;
wire   [0:0] icmp_ln1019_49_fu_6245_p2;
wire   [0:0] icmp_ln878_24_fu_6250_p2;
wire   [0:0] tmp_192_fu_6263_p3;
wire   [0:0] icmp_ln1019_48_fu_6240_p2;
wire   [0:0] xor_ln890_29_fu_6270_p2;
wire   [0:0] and_ln890_23_fu_6276_p2;
wire   [0:0] select_ln888_24_fu_6255_p3;
wire   [0:0] xor_ln895_53_fu_6296_p2;
wire   [0:0] or_ln895_23_fu_6302_p2;
wire   [0:0] xor_ln895_54_fu_6308_p2;
wire   [0:0] select_ln890_24_fu_6282_p3;
wire   [0:0] xor_ln896_63_fu_6319_p2;
wire   [0:0] and_ln891_23_fu_6290_p2;
wire   [0:0] or_ln896_23_fu_6325_p2;
wire   [0:0] xor_ln896_82_fu_6331_p2;
wire   [0:0] and_ln895_26_fu_6313_p2;
wire   [0:0] and_ln896_26_fu_6337_p2;
wire   [0:0] or_ln346_26_fu_6350_p2;
wire   [31:0] select_ln346_47_fu_6342_p3;
wire   [0:0] icmp_ln1420_1_fu_6369_p2;
wire   [0:0] icmp_ln1420_2_fu_6374_p2;
wire   [0:0] or_ln1420_fu_6379_p2;
wire   [0:0] icmp_ln1420_fu_6364_p2;
wire   [0:0] or_ln1420_1_fu_6385_p2;
wire   [31:0] temp1_V_3_9_fu_6356_p3;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter1_reg;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg    ap_loop_exit_ready_pp0_iter4_reg;
reg    ap_loop_exit_ready_pp0_iter5_reg;
reg    ap_loop_exit_ready_pp0_iter6_reg;
reg    ap_loop_exit_ready_pp0_iter7_reg;
reg    ap_loop_exit_ready_pp0_iter8_reg;
reg    ap_loop_exit_ready_pp0_iter9_reg;
reg    ap_loop_exit_ready_pp0_iter10_reg;
reg    ap_loop_exit_ready_pp0_iter11_reg;
reg    ap_loop_exit_ready_pp0_iter12_reg;
reg    ap_loop_exit_ready_pp0_iter13_reg;
reg    ap_loop_exit_ready_pp0_iter14_reg;
reg    ap_loop_exit_ready_pp0_iter15_reg;
reg    ap_loop_exit_ready_pp0_iter16_reg;
reg    ap_loop_exit_ready_pp0_iter17_reg;
reg    ap_loop_exit_ready_pp0_iter18_reg;
reg    ap_loop_exit_ready_pp0_iter19_reg;
reg    ap_loop_exit_ready_pp0_iter20_reg;
reg    ap_loop_exit_ready_pp0_iter21_reg;
reg    ap_loop_exit_ready_pp0_iter22_reg;
reg    ap_loop_exit_ready_pp0_iter23_reg;
reg    ap_loop_exit_ready_pp0_iter24_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
#0 ap_enable_reg_pp0_iter23 = 1'b0;
#0 ap_enable_reg_pp0_iter24 = 1'b0;
#0 ap_enable_reg_pp0_iter25 = 1'b0;
#0 ap_done_reg = 1'b0;
end

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U46(
    .din0(32'd4294938517),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_fu_526_p1),
    .dout(tmp_3_fu_530_p6)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U47(
    .din0(32'd4294966981),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_fu_526_p1),
    .dout(tmp_fu_544_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U48(
    .din0(mul_ln1273_fu_566_p0),
    .din1(tmp_3_reg_6651),
    .dout(mul_ln1273_fu_566_p2)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U49(
    .din0(mul_ln1273_1_fu_628_p0),
    .din1(tmp_reg_6656),
    .dout(mul_ln1273_1_fu_628_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U50(
    .din0(32'd4294951137),
    .din1(32'd4294938517),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622),
    .dout(tmp_6_fu_641_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U51(
    .din0(mul_ln1273_3_fu_871_p0),
    .din1(tmp_6_reg_6708),
    .dout(mul_ln1273_3_fu_871_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U52(
    .din0(32'd4294966543),
    .din1(32'd4294966981),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter1_reg),
    .dout(tmp_9_fu_884_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U53(
    .din0(mul_ln1273_6_fu_1114_p0),
    .din1(tmp_9_reg_6755),
    .dout(mul_ln1273_6_fu_1114_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U54(
    .din0(32'd4294958223),
    .din1(32'd4294951137),
    .din2(32'd4294938517),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter2_reg),
    .dout(tmp_s_fu_1127_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U55(
    .din0(mul_ln1273_7_fu_1357_p0),
    .din1(tmp_s_reg_6802),
    .dout(mul_ln1273_7_fu_1357_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U56(
    .din0(32'd4294966298),
    .din1(32'd4294966543),
    .din2(32'd4294966981),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter3_reg),
    .dout(tmp_14_fu_1370_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U57(
    .din0(mul_ln1273_8_fu_1600_p0),
    .din1(tmp_14_reg_6849),
    .dout(mul_ln1273_8_fu_1600_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U58(
    .din0(32'd4294962202),
    .din1(32'd4294958223),
    .din2(32'd4294951137),
    .din3(32'd4294938517),
    .din4(trunc_ln25_reg_6622_pp0_iter4_reg),
    .dout(tmp_17_fu_1613_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U59(
    .din0(mul_ln1273_9_fu_1843_p0),
    .din1(tmp_17_reg_6896),
    .dout(mul_ln1273_9_fu_1843_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U60(
    .din0(32'd4294966160),
    .din1(32'd4294966298),
    .din2(32'd4294966543),
    .din3(32'd4294966981),
    .din4(trunc_ln25_reg_6622_pp0_iter5_reg),
    .dout(tmp_20_fu_1856_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U61(
    .din0(mul_ln1273_10_fu_2086_p0),
    .din1(tmp_20_reg_6943),
    .dout(mul_ln1273_10_fu_2086_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U62(
    .din0(32'd28779),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter6_reg),
    .dout(tmp_23_fu_2099_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U63(
    .din0(mul_ln1273_11_fu_2329_p0),
    .din1(tmp_23_reg_6990),
    .dout(mul_ln1273_11_fu_2329_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U64(
    .din0(32'd315),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter7_reg),
    .dout(tmp_26_fu_2342_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U65(
    .din0(mul_ln1273_12_fu_2572_p0),
    .din1(tmp_26_reg_7037),
    .dout(mul_ln1273_12_fu_2572_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U66(
    .din0(32'd16159),
    .din1(32'd28779),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter8_reg),
    .dout(tmp_29_fu_2585_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U67(
    .din0(mul_ln1273_13_fu_2815_p0),
    .din1(tmp_29_reg_7084),
    .dout(mul_ln1273_13_fu_2815_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U68(
    .din0(32'd753),
    .din1(32'd315),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter9_reg),
    .dout(tmp_32_fu_2828_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U69(
    .din0(mul_ln1273_14_fu_3058_p0),
    .din1(tmp_32_reg_7131),
    .dout(mul_ln1273_14_fu_3058_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U70(
    .din0(32'd9073),
    .din1(32'd16159),
    .din2(32'd28779),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter10_reg),
    .dout(tmp_35_fu_3071_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U71(
    .din0(mul_ln1273_15_fu_3301_p0),
    .din1(tmp_35_reg_7178),
    .dout(mul_ln1273_15_fu_3301_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U72(
    .din0(32'd998),
    .din1(32'd753),
    .din2(32'd315),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter11_reg),
    .dout(tmp_38_fu_3314_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U73(
    .din0(mul_ln1273_16_fu_3544_p0),
    .din1(tmp_38_reg_7225),
    .dout(mul_ln1273_16_fu_3544_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U74(
    .din0(32'd5094),
    .din1(32'd9073),
    .din2(32'd16159),
    .din3(32'd28779),
    .din4(trunc_ln25_reg_6622_pp0_iter12_reg),
    .dout(tmp_41_fu_3557_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U75(
    .din0(mul_ln1273_17_fu_3787_p0),
    .din1(tmp_41_reg_7272),
    .dout(mul_ln1273_17_fu_3787_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U76(
    .din0(32'd1136),
    .din1(32'd998),
    .din2(32'd753),
    .din3(32'd315),
    .din4(trunc_ln25_reg_6622_pp0_iter13_reg),
    .dout(tmp_44_fu_3800_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U77(
    .din0(mul_ln1273_18_fu_4030_p0),
    .din1(tmp_44_reg_7319),
    .dout(mul_ln1273_18_fu_4030_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U78(
    .din0(32'd4294925214),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter14_reg),
    .dout(tmp_47_fu_4043_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U79(
    .din0(mul_ln1273_19_fu_4273_p0),
    .din1(tmp_47_reg_7366),
    .dout(mul_ln1273_19_fu_4273_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U80(
    .din0(32'd0),
    .din1(32'd4294925214),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter15_reg),
    .dout(tmp_50_fu_4286_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U81(
    .din0(mul_ln1273_20_fu_4516_p0),
    .din1(tmp_50_reg_7413),
    .dout(mul_ln1273_20_fu_4516_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U82(
    .din0(32'd0),
    .din1(32'd0),
    .din2(32'd4294925214),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter16_reg),
    .dout(tmp_53_fu_4529_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U83(
    .din0(mul_ln1273_21_fu_4759_p0),
    .din1(tmp_53_reg_7460),
    .dout(mul_ln1273_21_fu_4759_p2)
);

mpc_mux_42_32_1_1_x #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_x_U84(
    .din0(32'd0),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd4294925214),
    .din4(trunc_ln25_reg_6622_pp0_iter17_reg),
    .dout(tmp_56_fu_4772_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U85(
    .din0(mul_ln1273_22_fu_5002_p0),
    .din1(tmp_56_reg_7507),
    .dout(mul_ln1273_22_fu_5002_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U86(
    .din0(32'd42082),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter18_reg),
    .dout(tmp_59_fu_5015_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U87(
    .din0(mul_ln1273_23_fu_5245_p0),
    .din1(tmp_59_reg_7554),
    .dout(mul_ln1273_23_fu_5245_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U88(
    .din0(32'd0),
    .din1(32'd42082),
    .din2(32'd0),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter19_reg),
    .dout(tmp_62_fu_5258_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U89(
    .din0(mul_ln1273_24_fu_5488_p0),
    .din1(tmp_62_reg_7601),
    .dout(mul_ln1273_24_fu_5488_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U90(
    .din0(32'd0),
    .din1(32'd0),
    .din2(32'd42082),
    .din3(32'd0),
    .din4(trunc_ln25_reg_6622_pp0_iter20_reg),
    .dout(tmp_65_fu_5501_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U91(
    .din0(mul_ln1273_25_fu_5731_p0),
    .din1(tmp_65_reg_7648),
    .dout(mul_ln1273_25_fu_5731_p2)
);

mpc_mux_42_32_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .din2_WIDTH( 32 ),
    .din3_WIDTH( 32 ),
    .din4_WIDTH( 2 ),
    .dout_WIDTH( 32 ))
mux_42_32_1_1_U92(
    .din0(32'd0),
    .din1(32'd0),
    .din2(32'd0),
    .din3(32'd42082),
    .din4(trunc_ln25_reg_6622_pp0_iter21_reg),
    .dout(tmp_68_fu_5744_p6)
);

mpc_mul_32s_32s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 32 ),
    .dout_WIDTH( 64 ))
mul_32s_32s_64_1_1_U93(
    .din0(mul_ln1273_26_fu_5974_p0),
    .din1(tmp_68_reg_7695),
    .dout(mul_ln1273_26_fu_5974_p2)
);

mpc_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready_pp0_iter24_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter23 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter24 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter25 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln24_fu_514_p2 == 1'd0))) begin
            i_2_fu_174 <= add_ln24_fu_520_p2;
        end else if ((ap_loop_init == 1'b1)) begin
            i_2_fu_174 <= 3'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            temp1_V_3_1_fu_190 <= temp1_V_3_04;
        end else if ((ap_enable_reg_pp0_iter25 == 1'b1)) begin
            temp1_V_3_1_fu_190 <= temp1_V_3_fu_6391_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            temp1_V_3_2_fu_178 <= temp1_V_0_01;
        end else if ((ap_enable_reg_pp0_iter25 == 1'b1)) begin
            temp1_V_3_2_fu_178 <= temp1_V_3_8_fu_6415_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            temp1_V_3_3_fu_182 <= temp1_V_1_02;
        end else if ((ap_enable_reg_pp0_iter25 == 1'b1)) begin
            temp1_V_3_3_fu_182 <= temp1_V_3_7_fu_6407_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            temp1_V_3_4_fu_186 <= temp1_V_2_03;
        end else if ((ap_enable_reg_pp0_iter25 == 1'b1)) begin
            temp1_V_3_4_fu_186 <= temp1_V_3_6_fu_6399_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln1347_10_reg_7136 <= add_ln1347_10_fu_3004_p2;
        add_ln1347_11_reg_7183 <= add_ln1347_11_fu_3247_p2;
        add_ln1347_12_reg_7230 <= add_ln1347_12_fu_3490_p2;
        add_ln1347_13_reg_7277 <= add_ln1347_13_fu_3733_p2;
        add_ln1347_14_reg_7324 <= add_ln1347_14_fu_3976_p2;
        add_ln1347_15_reg_7371 <= add_ln1347_15_fu_4219_p2;
        add_ln1347_16_reg_7418 <= add_ln1347_16_fu_4462_p2;
        add_ln1347_17_reg_7465 <= add_ln1347_17_fu_4705_p2;
        add_ln1347_18_reg_7512 <= add_ln1347_18_fu_4948_p2;
        add_ln1347_19_reg_7559 <= add_ln1347_19_fu_5191_p2;
        add_ln1347_1_reg_6760 <= add_ln1347_1_fu_1060_p2;
        add_ln1347_20_reg_7606 <= add_ln1347_20_fu_5434_p2;
        add_ln1347_21_reg_7653 <= add_ln1347_21_fu_5677_p2;
        add_ln1347_22_reg_7700 <= add_ln1347_22_fu_5920_p2;
        add_ln1347_23_reg_7742 <= add_ln1347_23_fu_6150_p2;
        add_ln1347_3_reg_6807 <= add_ln1347_3_fu_1303_p2;
        add_ln1347_4_reg_6854 <= add_ln1347_4_fu_1546_p2;
        add_ln1347_5_reg_6901 <= add_ln1347_5_fu_1789_p2;
        add_ln1347_6_reg_6948 <= add_ln1347_6_fu_2032_p2;
        add_ln1347_7_reg_6995 <= add_ln1347_7_fu_2275_p2;
        add_ln1347_8_reg_7042 <= add_ln1347_8_fu_2518_p2;
        add_ln1347_9_reg_7089 <= add_ln1347_9_fu_2761_p2;
        add_ln1347_reg_6713 <= add_ln1347_fu_817_p2;
        ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
        ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
        ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
        ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
        ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
        ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
        ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
        ap_loop_exit_ready_pp0_iter17_reg <= ap_loop_exit_ready_pp0_iter16_reg;
        ap_loop_exit_ready_pp0_iter18_reg <= ap_loop_exit_ready_pp0_iter17_reg;
        ap_loop_exit_ready_pp0_iter19_reg <= ap_loop_exit_ready_pp0_iter18_reg;
        ap_loop_exit_ready_pp0_iter20_reg <= ap_loop_exit_ready_pp0_iter19_reg;
        ap_loop_exit_ready_pp0_iter21_reg <= ap_loop_exit_ready_pp0_iter20_reg;
        ap_loop_exit_ready_pp0_iter22_reg <= ap_loop_exit_ready_pp0_iter21_reg;
        ap_loop_exit_ready_pp0_iter23_reg <= ap_loop_exit_ready_pp0_iter22_reg;
        ap_loop_exit_ready_pp0_iter24_reg <= ap_loop_exit_ready_pp0_iter23_reg;
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        icmp_ln24_reg_6618_pp0_iter10_reg <= icmp_ln24_reg_6618_pp0_iter9_reg;
        icmp_ln24_reg_6618_pp0_iter11_reg <= icmp_ln24_reg_6618_pp0_iter10_reg;
        icmp_ln24_reg_6618_pp0_iter12_reg <= icmp_ln24_reg_6618_pp0_iter11_reg;
        icmp_ln24_reg_6618_pp0_iter13_reg <= icmp_ln24_reg_6618_pp0_iter12_reg;
        icmp_ln24_reg_6618_pp0_iter14_reg <= icmp_ln24_reg_6618_pp0_iter13_reg;
        icmp_ln24_reg_6618_pp0_iter15_reg <= icmp_ln24_reg_6618_pp0_iter14_reg;
        icmp_ln24_reg_6618_pp0_iter16_reg <= icmp_ln24_reg_6618_pp0_iter15_reg;
        icmp_ln24_reg_6618_pp0_iter17_reg <= icmp_ln24_reg_6618_pp0_iter16_reg;
        icmp_ln24_reg_6618_pp0_iter18_reg <= icmp_ln24_reg_6618_pp0_iter17_reg;
        icmp_ln24_reg_6618_pp0_iter19_reg <= icmp_ln24_reg_6618_pp0_iter18_reg;
        icmp_ln24_reg_6618_pp0_iter20_reg <= icmp_ln24_reg_6618_pp0_iter19_reg;
        icmp_ln24_reg_6618_pp0_iter21_reg <= icmp_ln24_reg_6618_pp0_iter20_reg;
        icmp_ln24_reg_6618_pp0_iter22_reg <= icmp_ln24_reg_6618_pp0_iter21_reg;
        icmp_ln24_reg_6618_pp0_iter23_reg <= icmp_ln24_reg_6618_pp0_iter22_reg;
        icmp_ln24_reg_6618_pp0_iter2_reg <= icmp_ln24_reg_6618_pp0_iter1_reg;
        icmp_ln24_reg_6618_pp0_iter3_reg <= icmp_ln24_reg_6618_pp0_iter2_reg;
        icmp_ln24_reg_6618_pp0_iter4_reg <= icmp_ln24_reg_6618_pp0_iter3_reg;
        icmp_ln24_reg_6618_pp0_iter5_reg <= icmp_ln24_reg_6618_pp0_iter4_reg;
        icmp_ln24_reg_6618_pp0_iter6_reg <= icmp_ln24_reg_6618_pp0_iter5_reg;
        icmp_ln24_reg_6618_pp0_iter7_reg <= icmp_ln24_reg_6618_pp0_iter6_reg;
        icmp_ln24_reg_6618_pp0_iter8_reg <= icmp_ln24_reg_6618_pp0_iter7_reg;
        icmp_ln24_reg_6618_pp0_iter9_reg <= icmp_ln24_reg_6618_pp0_iter8_reg;
        mul_ln1273_10_reg_6980 <= mul_ln1273_10_fu_2086_p2;
        mul_ln1273_11_reg_7027 <= mul_ln1273_11_fu_2329_p2;
        mul_ln1273_12_reg_7074 <= mul_ln1273_12_fu_2572_p2;
        mul_ln1273_13_reg_7121 <= mul_ln1273_13_fu_2815_p2;
        mul_ln1273_14_reg_7168 <= mul_ln1273_14_fu_3058_p2;
        mul_ln1273_15_reg_7215 <= mul_ln1273_15_fu_3301_p2;
        mul_ln1273_16_reg_7262 <= mul_ln1273_16_fu_3544_p2;
        mul_ln1273_17_reg_7309 <= mul_ln1273_17_fu_3787_p2;
        mul_ln1273_18_reg_7356 <= mul_ln1273_18_fu_4030_p2;
        mul_ln1273_19_reg_7403 <= mul_ln1273_19_fu_4273_p2;
        mul_ln1273_20_reg_7450 <= mul_ln1273_20_fu_4516_p2;
        mul_ln1273_21_reg_7497 <= mul_ln1273_21_fu_4759_p2;
        mul_ln1273_22_reg_7544 <= mul_ln1273_22_fu_5002_p2;
        mul_ln1273_23_reg_7591 <= mul_ln1273_23_fu_5245_p2;
        mul_ln1273_24_reg_7638 <= mul_ln1273_24_fu_5488_p2;
        mul_ln1273_25_reg_7685 <= mul_ln1273_25_fu_5731_p2;
        mul_ln1273_26_reg_7732 <= mul_ln1273_26_fu_5974_p2;
        mul_ln1273_3_reg_6745 <= mul_ln1273_3_fu_871_p2;
        mul_ln1273_6_reg_6792 <= mul_ln1273_6_fu_1114_p2;
        mul_ln1273_7_reg_6839 <= mul_ln1273_7_fu_1357_p2;
        mul_ln1273_8_reg_6886 <= mul_ln1273_8_fu_1600_p2;
        mul_ln1273_9_reg_6933 <= mul_ln1273_9_fu_1843_p2;
        tmp_100_reg_6891 <= mul_ln1273_8_fu_1600_p2[32'd15];
        tmp_100_reg_6891_pp0_iter6_reg <= tmp_100_reg_6891;
        tmp_103_reg_6953 <= add_ln1347_6_fu_2032_p2[32'd63];
        tmp_104_reg_6964 <= add_ln1347_6_fu_2032_p2[32'd47];
        tmp_105_reg_6938 <= mul_ln1273_9_fu_1843_p2[32'd15];
        tmp_105_reg_6938_pp0_iter7_reg <= tmp_105_reg_6938;
        tmp_108_reg_7000 <= add_ln1347_7_fu_2275_p2[32'd63];
        tmp_109_reg_7011 <= add_ln1347_7_fu_2275_p2[32'd47];
        tmp_10_reg_6828 <= {{add_ln1347_3_fu_1303_p2[63:49]}};
        tmp_110_reg_6985 <= mul_ln1273_10_fu_2086_p2[32'd15];
        tmp_110_reg_6985_pp0_iter8_reg <= tmp_110_reg_6985;
        tmp_113_reg_7047 <= add_ln1347_8_fu_2518_p2[32'd63];
        tmp_114_reg_7058 <= add_ln1347_8_fu_2518_p2[32'd47];
        tmp_115_reg_7032 <= mul_ln1273_11_fu_2329_p2[32'd15];
        tmp_115_reg_7032_pp0_iter9_reg <= tmp_115_reg_7032;
        tmp_118_reg_7094 <= add_ln1347_9_fu_2761_p2[32'd63];
        tmp_119_reg_7105 <= add_ln1347_9_fu_2761_p2[32'd47];
        tmp_11_reg_6833 <= {{add_ln1347_3_fu_1303_p2[63:48]}};
        tmp_120_reg_7079 <= mul_ln1273_12_fu_2572_p2[32'd15];
        tmp_120_reg_7079_pp0_iter10_reg <= tmp_120_reg_7079;
        tmp_123_reg_7141 <= add_ln1347_10_fu_3004_p2[32'd63];
        tmp_124_reg_7152 <= add_ln1347_10_fu_3004_p2[32'd47];
        tmp_125_reg_7126 <= mul_ln1273_13_fu_2815_p2[32'd15];
        tmp_125_reg_7126_pp0_iter11_reg <= tmp_125_reg_7126;
        tmp_128_reg_7188 <= add_ln1347_11_fu_3247_p2[32'd63];
        tmp_129_reg_7199 <= add_ln1347_11_fu_3247_p2[32'd47];
        tmp_12_reg_6875 <= {{add_ln1347_4_fu_1546_p2[63:49]}};
        tmp_130_reg_7173 <= mul_ln1273_14_fu_3058_p2[32'd15];
        tmp_130_reg_7173_pp0_iter12_reg <= tmp_130_reg_7173;
        tmp_133_reg_7235 <= add_ln1347_12_fu_3490_p2[32'd63];
        tmp_134_reg_7246 <= add_ln1347_12_fu_3490_p2[32'd47];
        tmp_135_reg_7220 <= mul_ln1273_15_fu_3301_p2[32'd15];
        tmp_135_reg_7220_pp0_iter13_reg <= tmp_135_reg_7220;
        tmp_138_reg_7282 <= add_ln1347_13_fu_3733_p2[32'd63];
        tmp_139_reg_7293 <= add_ln1347_13_fu_3733_p2[32'd47];
        tmp_13_reg_6880 <= {{add_ln1347_4_fu_1546_p2[63:48]}};
        tmp_140_reg_7267 <= mul_ln1273_16_fu_3544_p2[32'd15];
        tmp_140_reg_7267_pp0_iter14_reg <= tmp_140_reg_7267;
        tmp_143_reg_7329 <= add_ln1347_14_fu_3976_p2[32'd63];
        tmp_144_reg_7340 <= add_ln1347_14_fu_3976_p2[32'd47];
        tmp_145_reg_7314 <= mul_ln1273_17_fu_3787_p2[32'd15];
        tmp_145_reg_7314_pp0_iter15_reg <= tmp_145_reg_7314;
        tmp_148_reg_7376 <= add_ln1347_15_fu_4219_p2[32'd63];
        tmp_149_reg_7387 <= add_ln1347_15_fu_4219_p2[32'd47];
        tmp_14_reg_6849 <= tmp_14_fu_1370_p6;
        tmp_150_reg_7361 <= mul_ln1273_18_fu_4030_p2[32'd15];
        tmp_150_reg_7361_pp0_iter16_reg <= tmp_150_reg_7361;
        tmp_153_reg_7423 <= add_ln1347_16_fu_4462_p2[32'd63];
        tmp_154_reg_7434 <= add_ln1347_16_fu_4462_p2[32'd47];
        tmp_155_reg_7408 <= mul_ln1273_19_fu_4273_p2[32'd15];
        tmp_155_reg_7408_pp0_iter17_reg <= tmp_155_reg_7408;
        tmp_158_reg_7470 <= add_ln1347_17_fu_4705_p2[32'd63];
        tmp_159_reg_7481 <= add_ln1347_17_fu_4705_p2[32'd47];
        tmp_15_reg_6922 <= {{add_ln1347_5_fu_1789_p2[63:49]}};
        tmp_160_reg_7455 <= mul_ln1273_20_fu_4516_p2[32'd15];
        tmp_160_reg_7455_pp0_iter18_reg <= tmp_160_reg_7455;
        tmp_163_reg_7517 <= add_ln1347_18_fu_4948_p2[32'd63];
        tmp_164_reg_7528 <= add_ln1347_18_fu_4948_p2[32'd47];
        tmp_165_reg_7502 <= mul_ln1273_21_fu_4759_p2[32'd15];
        tmp_165_reg_7502_pp0_iter19_reg <= tmp_165_reg_7502;
        tmp_168_reg_7564 <= add_ln1347_19_fu_5191_p2[32'd63];
        tmp_169_reg_7575 <= add_ln1347_19_fu_5191_p2[32'd47];
        tmp_16_reg_6927 <= {{add_ln1347_5_fu_1789_p2[63:48]}};
        tmp_170_reg_7549 <= mul_ln1273_22_fu_5002_p2[32'd15];
        tmp_170_reg_7549_pp0_iter20_reg <= tmp_170_reg_7549;
        tmp_173_reg_7611 <= add_ln1347_20_fu_5434_p2[32'd63];
        tmp_174_reg_7622 <= add_ln1347_20_fu_5434_p2[32'd47];
        tmp_175_reg_7596 <= mul_ln1273_23_fu_5245_p2[32'd15];
        tmp_175_reg_7596_pp0_iter21_reg <= tmp_175_reg_7596;
        tmp_178_reg_7658 <= add_ln1347_21_fu_5677_p2[32'd63];
        tmp_179_reg_7669 <= add_ln1347_21_fu_5677_p2[32'd47];
        tmp_17_reg_6896 <= tmp_17_fu_1613_p6;
        tmp_180_reg_7643 <= mul_ln1273_24_fu_5488_p2[32'd15];
        tmp_180_reg_7643_pp0_iter22_reg <= tmp_180_reg_7643;
        tmp_183_reg_7705 <= add_ln1347_22_fu_5920_p2[32'd63];
        tmp_184_reg_7716 <= add_ln1347_22_fu_5920_p2[32'd47];
        tmp_185_reg_7690 <= mul_ln1273_25_fu_5731_p2[32'd15];
        tmp_185_reg_7690_pp0_iter23_reg <= tmp_185_reg_7690;
        tmp_188_reg_7747 <= add_ln1347_23_fu_6150_p2[32'd63];
        tmp_189_reg_7758 <= add_ln1347_23_fu_6150_p2[32'd47];
        tmp_18_reg_6969 <= {{add_ln1347_6_fu_2032_p2[63:49]}};
        tmp_190_reg_7737 <= mul_ln1273_26_fu_5974_p2[32'd15];
        tmp_190_reg_7737_pp0_iter24_reg <= tmp_190_reg_7737;
        tmp_19_reg_6974 <= {{add_ln1347_6_fu_2032_p2[63:48]}};
        tmp_20_reg_6943 <= tmp_20_fu_1856_p6;
        tmp_21_reg_7016 <= {{add_ln1347_7_fu_2275_p2[63:49]}};
        tmp_22_reg_7021 <= {{add_ln1347_7_fu_2275_p2[63:48]}};
        tmp_23_reg_6990 <= tmp_23_fu_2099_p6;
        tmp_24_reg_7063 <= {{add_ln1347_8_fu_2518_p2[63:49]}};
        tmp_25_reg_7068 <= {{add_ln1347_8_fu_2518_p2[63:48]}};
        tmp_26_reg_7037 <= tmp_26_fu_2342_p6;
        tmp_27_reg_7110 <= {{add_ln1347_9_fu_2761_p2[63:49]}};
        tmp_28_reg_7115 <= {{add_ln1347_9_fu_2761_p2[63:48]}};
        tmp_29_reg_7084 <= tmp_29_fu_2585_p6;
        tmp_30_reg_7157 <= {{add_ln1347_10_fu_3004_p2[63:49]}};
        tmp_31_reg_7162 <= {{add_ln1347_10_fu_3004_p2[63:48]}};
        tmp_32_reg_7131 <= tmp_32_fu_2828_p6;
        tmp_33_reg_7204 <= {{add_ln1347_11_fu_3247_p2[63:49]}};
        tmp_34_reg_7209 <= {{add_ln1347_11_fu_3247_p2[63:48]}};
        tmp_35_reg_7178 <= tmp_35_fu_3071_p6;
        tmp_36_reg_7251 <= {{add_ln1347_12_fu_3490_p2[63:49]}};
        tmp_37_reg_7256 <= {{add_ln1347_12_fu_3490_p2[63:48]}};
        tmp_38_reg_7225 <= tmp_38_fu_3314_p6;
        tmp_39_reg_7298 <= {{add_ln1347_13_fu_3733_p2[63:49]}};
        tmp_40_reg_7303 <= {{add_ln1347_13_fu_3733_p2[63:48]}};
        tmp_41_reg_7272 <= tmp_41_fu_3557_p6;
        tmp_42_reg_7345 <= {{add_ln1347_14_fu_3976_p2[63:49]}};
        tmp_43_reg_7350 <= {{add_ln1347_14_fu_3976_p2[63:48]}};
        tmp_44_reg_7319 <= tmp_44_fu_3800_p6;
        tmp_45_reg_7392 <= {{add_ln1347_15_fu_4219_p2[63:49]}};
        tmp_46_reg_7397 <= {{add_ln1347_15_fu_4219_p2[63:48]}};
        tmp_47_reg_7366 <= tmp_47_fu_4043_p6;
        tmp_48_reg_7439 <= {{add_ln1347_16_fu_4462_p2[63:49]}};
        tmp_49_reg_7444 <= {{add_ln1347_16_fu_4462_p2[63:48]}};
        tmp_4_reg_6734 <= {{add_ln1347_fu_817_p2[63:49]}};
        tmp_50_reg_7413 <= tmp_50_fu_4286_p6;
        tmp_51_reg_7486 <= {{add_ln1347_17_fu_4705_p2[63:49]}};
        tmp_52_reg_7491 <= {{add_ln1347_17_fu_4705_p2[63:48]}};
        tmp_53_reg_7460 <= tmp_53_fu_4529_p6;
        tmp_54_reg_7533 <= {{add_ln1347_18_fu_4948_p2[63:49]}};
        tmp_55_reg_7538 <= {{add_ln1347_18_fu_4948_p2[63:48]}};
        tmp_56_reg_7507 <= tmp_56_fu_4772_p6;
        tmp_57_reg_7580 <= {{add_ln1347_19_fu_5191_p2[63:49]}};
        tmp_58_reg_7585 <= {{add_ln1347_19_fu_5191_p2[63:48]}};
        tmp_59_reg_7554 <= tmp_59_fu_5015_p6;
        tmp_5_reg_6739 <= {{add_ln1347_fu_817_p2[63:48]}};
        tmp_60_reg_7627 <= {{add_ln1347_20_fu_5434_p2[63:49]}};
        tmp_61_reg_7632 <= {{add_ln1347_20_fu_5434_p2[63:48]}};
        tmp_62_reg_7601 <= tmp_62_fu_5258_p6;
        tmp_63_reg_7674 <= {{add_ln1347_21_fu_5677_p2[63:49]}};
        tmp_64_reg_7679 <= {{add_ln1347_21_fu_5677_p2[63:48]}};
        tmp_65_reg_7648 <= tmp_65_fu_5501_p6;
        tmp_66_reg_7721 <= {{add_ln1347_22_fu_5920_p2[63:49]}};
        tmp_67_reg_7726 <= {{add_ln1347_22_fu_5920_p2[63:48]}};
        tmp_68_reg_7695 <= tmp_68_fu_5744_p6;
        tmp_69_reg_7763 <= {{add_ln1347_23_fu_6150_p2[63:49]}};
        tmp_70_reg_7768 <= {{add_ln1347_23_fu_6150_p2[63:48]}};
        tmp_78_reg_6718 <= add_ln1347_fu_817_p2[32'd63];
        tmp_79_reg_6729 <= add_ln1347_fu_817_p2[32'd47];
        tmp_7_reg_6781 <= {{add_ln1347_1_fu_1060_p2[63:49]}};
        tmp_80_reg_6703_pp0_iter2_reg <= tmp_80_reg_6703;
        tmp_83_reg_6765 <= add_ln1347_1_fu_1060_p2[32'd63];
        tmp_84_reg_6776 <= add_ln1347_1_fu_1060_p2[32'd47];
        tmp_85_reg_6750 <= mul_ln1273_3_fu_871_p2[32'd15];
        tmp_85_reg_6750_pp0_iter3_reg <= tmp_85_reg_6750;
        tmp_88_reg_6812 <= add_ln1347_3_fu_1303_p2[32'd63];
        tmp_89_reg_6823 <= add_ln1347_3_fu_1303_p2[32'd47];
        tmp_8_reg_6786 <= {{add_ln1347_1_fu_1060_p2[63:48]}};
        tmp_90_reg_6797 <= mul_ln1273_6_fu_1114_p2[32'd15];
        tmp_90_reg_6797_pp0_iter4_reg <= tmp_90_reg_6797;
        tmp_93_reg_6859 <= add_ln1347_4_fu_1546_p2[32'd63];
        tmp_94_reg_6870 <= add_ln1347_4_fu_1546_p2[32'd47];
        tmp_95_reg_6844 <= mul_ln1273_7_fu_1357_p2[32'd15];
        tmp_95_reg_6844_pp0_iter5_reg <= tmp_95_reg_6844;
        tmp_98_reg_6906 <= add_ln1347_5_fu_1789_p2[32'd63];
        tmp_99_reg_6917 <= add_ln1347_5_fu_1789_p2[32'd47];
        tmp_9_reg_6755 <= tmp_9_fu_884_p6;
        tmp_s_reg_6802 <= tmp_s_fu_1127_p6;
        trunc_ln25_reg_6622_pp0_iter10_reg <= trunc_ln25_reg_6622_pp0_iter9_reg;
        trunc_ln25_reg_6622_pp0_iter11_reg <= trunc_ln25_reg_6622_pp0_iter10_reg;
        trunc_ln25_reg_6622_pp0_iter12_reg <= trunc_ln25_reg_6622_pp0_iter11_reg;
        trunc_ln25_reg_6622_pp0_iter13_reg <= trunc_ln25_reg_6622_pp0_iter12_reg;
        trunc_ln25_reg_6622_pp0_iter14_reg <= trunc_ln25_reg_6622_pp0_iter13_reg;
        trunc_ln25_reg_6622_pp0_iter15_reg <= trunc_ln25_reg_6622_pp0_iter14_reg;
        trunc_ln25_reg_6622_pp0_iter16_reg <= trunc_ln25_reg_6622_pp0_iter15_reg;
        trunc_ln25_reg_6622_pp0_iter17_reg <= trunc_ln25_reg_6622_pp0_iter16_reg;
        trunc_ln25_reg_6622_pp0_iter18_reg <= trunc_ln25_reg_6622_pp0_iter17_reg;
        trunc_ln25_reg_6622_pp0_iter19_reg <= trunc_ln25_reg_6622_pp0_iter18_reg;
        trunc_ln25_reg_6622_pp0_iter20_reg <= trunc_ln25_reg_6622_pp0_iter19_reg;
        trunc_ln25_reg_6622_pp0_iter21_reg <= trunc_ln25_reg_6622_pp0_iter20_reg;
        trunc_ln25_reg_6622_pp0_iter22_reg <= trunc_ln25_reg_6622_pp0_iter21_reg;
        trunc_ln25_reg_6622_pp0_iter23_reg <= trunc_ln25_reg_6622_pp0_iter22_reg;
        trunc_ln25_reg_6622_pp0_iter24_reg <= trunc_ln25_reg_6622_pp0_iter23_reg;
        trunc_ln25_reg_6622_pp0_iter2_reg <= trunc_ln25_reg_6622_pp0_iter1_reg;
        trunc_ln25_reg_6622_pp0_iter3_reg <= trunc_ln25_reg_6622_pp0_iter2_reg;
        trunc_ln25_reg_6622_pp0_iter4_reg <= trunc_ln25_reg_6622_pp0_iter3_reg;
        trunc_ln25_reg_6622_pp0_iter5_reg <= trunc_ln25_reg_6622_pp0_iter4_reg;
        trunc_ln25_reg_6622_pp0_iter6_reg <= trunc_ln25_reg_6622_pp0_iter5_reg;
        trunc_ln25_reg_6622_pp0_iter7_reg <= trunc_ln25_reg_6622_pp0_iter6_reg;
        trunc_ln25_reg_6622_pp0_iter8_reg <= trunc_ln25_reg_6622_pp0_iter7_reg;
        trunc_ln25_reg_6622_pp0_iter9_reg <= trunc_ln25_reg_6622_pp0_iter8_reg;
        trunc_ln818_10_reg_7194 <= {{add_ln1347_11_fu_3247_p2[47:16]}};
        trunc_ln818_11_reg_7241 <= {{add_ln1347_12_fu_3490_p2[47:16]}};
        trunc_ln818_12_reg_7288 <= {{add_ln1347_13_fu_3733_p2[47:16]}};
        trunc_ln818_13_reg_7335 <= {{add_ln1347_14_fu_3976_p2[47:16]}};
        trunc_ln818_14_reg_7382 <= {{add_ln1347_15_fu_4219_p2[47:16]}};
        trunc_ln818_15_reg_7429 <= {{add_ln1347_16_fu_4462_p2[47:16]}};
        trunc_ln818_16_reg_7476 <= {{add_ln1347_17_fu_4705_p2[47:16]}};
        trunc_ln818_17_reg_7523 <= {{add_ln1347_18_fu_4948_p2[47:16]}};
        trunc_ln818_18_reg_7570 <= {{add_ln1347_19_fu_5191_p2[47:16]}};
        trunc_ln818_19_reg_7617 <= {{add_ln1347_20_fu_5434_p2[47:16]}};
        trunc_ln818_1_reg_6724 <= {{add_ln1347_fu_817_p2[47:16]}};
        trunc_ln818_20_reg_7664 <= {{add_ln1347_21_fu_5677_p2[47:16]}};
        trunc_ln818_21_reg_7711 <= {{add_ln1347_22_fu_5920_p2[47:16]}};
        trunc_ln818_22_reg_7753 <= {{add_ln1347_23_fu_6150_p2[47:16]}};
        trunc_ln818_2_reg_6959 <= {{add_ln1347_6_fu_2032_p2[47:16]}};
        trunc_ln818_3_reg_6771 <= {{add_ln1347_1_fu_1060_p2[47:16]}};
        trunc_ln818_4_reg_7006 <= {{add_ln1347_7_fu_2275_p2[47:16]}};
        trunc_ln818_5_reg_7053 <= {{add_ln1347_8_fu_2518_p2[47:16]}};
        trunc_ln818_6_reg_6818 <= {{add_ln1347_3_fu_1303_p2[47:16]}};
        trunc_ln818_7_reg_7100 <= {{add_ln1347_9_fu_2761_p2[47:16]}};
        trunc_ln818_8_reg_7147 <= {{add_ln1347_10_fu_3004_p2[47:16]}};
        trunc_ln818_9_reg_6865 <= {{add_ln1347_4_fu_1546_p2[47:16]}};
        trunc_ln818_s_reg_6912 <= {{add_ln1347_5_fu_1789_p2[47:16]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        icmp_ln24_reg_6618 <= icmp_ln24_fu_514_p2;
        icmp_ln24_reg_6618_pp0_iter1_reg <= icmp_ln24_reg_6618;
        mul_ln1273_1_reg_6698 <= mul_ln1273_1_fu_628_p2;
        mul_ln1273_reg_6661 <= mul_ln1273_fu_566_p2;
        sext_ln1273_10_cast_reg_6563 <= sext_ln1273_10_cast_fu_442_p1;
        sext_ln1273_11_cast_reg_6558 <= sext_ln1273_11_cast_fu_438_p1;
        sext_ln1273_12_cast_reg_6553 <= sext_ln1273_12_cast_fu_434_p1;
        sext_ln1273_13_cast_reg_6548 <= sext_ln1273_13_cast_fu_430_p1;
        sext_ln1273_14_cast_reg_6543 <= sext_ln1273_14_cast_fu_426_p1;
        sext_ln1273_15_cast_reg_6538 <= sext_ln1273_15_cast_fu_422_p1;
        sext_ln1273_16_cast_reg_6533 <= sext_ln1273_16_cast_fu_418_p1;
        sext_ln1273_17_cast_reg_6528 <= sext_ln1273_17_cast_fu_414_p1;
        sext_ln1273_18_cast_reg_6523 <= sext_ln1273_18_cast_fu_410_p1;
        sext_ln1273_19_cast_reg_6518 <= sext_ln1273_19_cast_fu_406_p1;
        sext_ln1273_1_cast_reg_6608 <= sext_ln1273_1_cast_fu_478_p1;
        sext_ln1273_20_cast_reg_6513 <= sext_ln1273_20_cast_fu_402_p1;
        sext_ln1273_21_cast_reg_6508 <= sext_ln1273_21_cast_fu_398_p1;
        sext_ln1273_22_cast_reg_6503 <= sext_ln1273_22_cast_fu_394_p1;
        sext_ln1273_23_cast_reg_6498 <= sext_ln1273_23_cast_fu_390_p1;
        sext_ln1273_24_cast_reg_6603 <= sext_ln1273_24_cast_fu_474_p1;
        sext_ln1273_3_cast_reg_6598 <= sext_ln1273_3_cast_fu_470_p1;
        sext_ln1273_4_cast_reg_6593 <= sext_ln1273_4_cast_fu_466_p1;
        sext_ln1273_5_cast_reg_6588 <= sext_ln1273_5_cast_fu_462_p1;
        sext_ln1273_6_cast_reg_6583 <= sext_ln1273_6_cast_fu_458_p1;
        sext_ln1273_7_cast_reg_6578 <= sext_ln1273_7_cast_fu_454_p1;
        sext_ln1273_8_cast_reg_6573 <= sext_ln1273_8_cast_fu_450_p1;
        sext_ln1273_9_cast_reg_6568 <= sext_ln1273_9_cast_fu_446_p1;
        sext_ln1273_cast_reg_6613 <= sext_ln1273_cast_fu_482_p1;
        tmp_1_reg_6687 <= {{mul_ln1273_fu_566_p2[63:49]}};
        tmp_2_reg_6692 <= {{mul_ln1273_fu_566_p2[63:48]}};
        tmp_6_reg_6708 <= tmp_6_fu_641_p6;
        tmp_73_reg_6666 <= mul_ln1273_fu_566_p2[32'd63];
        tmp_74_reg_6677 <= mul_ln1273_fu_566_p2[32'd47];
        tmp_75_reg_6682 <= mul_ln1273_fu_566_p2[32'd15];
        tmp_80_reg_6703 <= mul_ln1273_1_fu_628_p2[32'd15];
        trunc_ln1_reg_6672 <= {{mul_ln1273_fu_566_p2[47:16]}};
        trunc_ln25_reg_6622_pp0_iter1_reg <= trunc_ln25_reg_6622;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln24_fu_514_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_3_reg_6651 <= tmp_3_fu_530_p6;
        tmp_reg_6656 <= tmp_fu_544_p6;
        trunc_ln25_reg_6622 <= trunc_ln25_fu_526_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln24_fu_514_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_condition_exit_pp0_iter0_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter0_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready_pp0_iter24_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0) & (ap_loop_init == 1'b1))) begin
        ap_sig_allocacmp_i = 3'd0;
    end else begin
        ap_sig_allocacmp_i = i_2_fu_174;
    end
end

always @ (*) begin
    if (((icmp_ln24_reg_6618_pp0_iter23_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        temp1_V_0_1_out_ap_vld = 1'b1;
    end else begin
        temp1_V_0_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln24_reg_6618_pp0_iter23_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        temp1_V_1_1_out_ap_vld = 1'b1;
    end else begin
        temp1_V_1_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln24_reg_6618_pp0_iter23_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        temp1_V_2_1_out_ap_vld = 1'b1;
    end else begin
        temp1_V_2_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln24_reg_6618_pp0_iter23_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        temp1_V_3_1_out_ap_vld = 1'b1;
    end else begin
        temp1_V_3_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln1347_10_fu_3004_p2 = ($signed(sext_ln813_11_fu_3000_p1) + $signed(mul_ln1273_13_reg_7121));

assign add_ln1347_11_fu_3247_p2 = ($signed(sext_ln813_12_fu_3243_p1) + $signed(mul_ln1273_14_reg_7168));

assign add_ln1347_12_fu_3490_p2 = ($signed(sext_ln813_13_fu_3486_p1) + $signed(mul_ln1273_15_reg_7215));

assign add_ln1347_13_fu_3733_p2 = ($signed(sext_ln813_14_fu_3729_p1) + $signed(mul_ln1273_16_reg_7262));

assign add_ln1347_14_fu_3976_p2 = ($signed(sext_ln813_15_fu_3972_p1) + $signed(mul_ln1273_17_reg_7309));

assign add_ln1347_15_fu_4219_p2 = ($signed(sext_ln813_16_fu_4215_p1) + $signed(mul_ln1273_18_reg_7356));

assign add_ln1347_16_fu_4462_p2 = ($signed(sext_ln813_17_fu_4458_p1) + $signed(mul_ln1273_19_reg_7403));

assign add_ln1347_17_fu_4705_p2 = ($signed(sext_ln813_18_fu_4701_p1) + $signed(mul_ln1273_20_reg_7450));

assign add_ln1347_18_fu_4948_p2 = ($signed(sext_ln813_19_fu_4944_p1) + $signed(mul_ln1273_21_reg_7497));

assign add_ln1347_19_fu_5191_p2 = ($signed(sext_ln813_20_fu_5187_p1) + $signed(mul_ln1273_22_reg_7544));

assign add_ln1347_1_fu_1060_p2 = ($signed(sext_ln813_4_fu_1056_p1) + $signed(mul_ln1273_3_reg_6745));

assign add_ln1347_20_fu_5434_p2 = ($signed(sext_ln813_21_fu_5430_p1) + $signed(mul_ln1273_23_reg_7591));

assign add_ln1347_21_fu_5677_p2 = ($signed(sext_ln813_22_fu_5673_p1) + $signed(mul_ln1273_24_reg_7638));

assign add_ln1347_22_fu_5920_p2 = ($signed(sext_ln813_23_fu_5916_p1) + $signed(mul_ln1273_25_reg_7685));

assign add_ln1347_23_fu_6150_p2 = ($signed(sext_ln813_24_fu_6146_p1) + $signed(mul_ln1273_26_reg_7732));

assign add_ln1347_3_fu_1303_p2 = ($signed(sext_ln813_5_fu_1299_p1) + $signed(mul_ln1273_6_reg_6792));

assign add_ln1347_4_fu_1546_p2 = ($signed(sext_ln813_6_fu_1542_p1) + $signed(mul_ln1273_7_reg_6839));

assign add_ln1347_5_fu_1789_p2 = ($signed(sext_ln813_7_fu_1785_p1) + $signed(mul_ln1273_8_reg_6886));

assign add_ln1347_6_fu_2032_p2 = ($signed(sext_ln813_8_fu_2028_p1) + $signed(mul_ln1273_9_reg_6933));

assign add_ln1347_7_fu_2275_p2 = ($signed(sext_ln813_fu_2271_p1) + $signed(mul_ln1273_10_reg_6980));

assign add_ln1347_8_fu_2518_p2 = ($signed(sext_ln813_9_fu_2514_p1) + $signed(mul_ln1273_11_reg_7027));

assign add_ln1347_9_fu_2761_p2 = ($signed(sext_ln813_10_fu_2757_p1) + $signed(mul_ln1273_12_reg_7074));

assign add_ln1347_fu_817_p2 = ($signed(sext_ln813_3_fu_813_p1) + $signed(mul_ln1273_1_reg_6698));

assign add_ln24_fu_520_p2 = (ap_sig_allocacmp_i + 3'd1);

assign add_ln377_10_fu_2358_p2 = (zext_ln377_7_fu_2355_p1 + trunc_ln818_4_reg_7006);

assign add_ln377_11_fu_2601_p2 = (zext_ln377_8_fu_2598_p1 + trunc_ln818_5_reg_7053);

assign add_ln377_12_fu_2844_p2 = (zext_ln377_9_fu_2841_p1 + trunc_ln818_7_reg_7100);

assign add_ln377_13_fu_3087_p2 = (zext_ln377_10_fu_3084_p1 + trunc_ln818_8_reg_7147);

assign add_ln377_14_fu_3330_p2 = (zext_ln377_11_fu_3327_p1 + trunc_ln818_10_reg_7194);

assign add_ln377_15_fu_3573_p2 = (zext_ln377_12_fu_3570_p1 + trunc_ln818_11_reg_7241);

assign add_ln377_16_fu_3816_p2 = (zext_ln377_13_fu_3813_p1 + trunc_ln818_12_reg_7288);

assign add_ln377_17_fu_4059_p2 = (zext_ln377_14_fu_4056_p1 + trunc_ln818_13_reg_7335);

assign add_ln377_18_fu_4302_p2 = (zext_ln377_15_fu_4299_p1 + trunc_ln818_14_reg_7382);

assign add_ln377_19_fu_4545_p2 = (zext_ln377_16_fu_4542_p1 + trunc_ln818_15_reg_7429);

assign add_ln377_1_fu_900_p2 = (zext_ln377_1_fu_897_p1 + trunc_ln818_1_reg_6724);

assign add_ln377_20_fu_4788_p2 = (zext_ln377_17_fu_4785_p1 + trunc_ln818_16_reg_7476);

assign add_ln377_21_fu_5031_p2 = (zext_ln377_18_fu_5028_p1 + trunc_ln818_17_reg_7523);

assign add_ln377_22_fu_5274_p2 = (zext_ln377_19_fu_5271_p1 + trunc_ln818_18_reg_7570);

assign add_ln377_23_fu_5517_p2 = (zext_ln377_20_fu_5514_p1 + trunc_ln818_19_reg_7617);

assign add_ln377_24_fu_5760_p2 = (zext_ln377_21_fu_5757_p1 + trunc_ln818_20_reg_7664);

assign add_ln377_25_fu_5990_p2 = (zext_ln377_22_fu_5987_p1 + trunc_ln818_21_reg_7711);

assign add_ln377_26_fu_6216_p2 = (zext_ln377_23_fu_6213_p1 + trunc_ln818_22_reg_7753);

assign add_ln377_3_fu_1143_p2 = (zext_ln377_2_fu_1140_p1 + trunc_ln818_3_reg_6771);

assign add_ln377_6_fu_1386_p2 = (zext_ln377_3_fu_1383_p1 + trunc_ln818_6_reg_6818);

assign add_ln377_7_fu_1629_p2 = (zext_ln377_4_fu_1626_p1 + trunc_ln818_9_reg_6865);

assign add_ln377_8_fu_1872_p2 = (zext_ln377_5_fu_1869_p1 + trunc_ln818_s_reg_6912);

assign add_ln377_9_fu_2115_p2 = (zext_ln377_6_fu_2112_p1 + trunc_ln818_2_reg_6959);

assign add_ln377_fu_657_p2 = (zext_ln377_fu_654_p1 + trunc_ln1_reg_6672);

assign and_ln378_10_fu_2377_p2 = (xor_ln896_30_fu_2371_p2 & tmp_109_reg_7011);

assign and_ln378_11_fu_2620_p2 = (xor_ln896_32_fu_2614_p2 & tmp_114_reg_7058);

assign and_ln378_12_fu_2863_p2 = (xor_ln896_34_fu_2857_p2 & tmp_119_reg_7105);

assign and_ln378_13_fu_3106_p2 = (xor_ln896_36_fu_3100_p2 & tmp_124_reg_7152);

assign and_ln378_14_fu_3349_p2 = (xor_ln896_38_fu_3343_p2 & tmp_129_reg_7199);

assign and_ln378_15_fu_3592_p2 = (xor_ln896_40_fu_3586_p2 & tmp_134_reg_7246);

assign and_ln378_16_fu_3835_p2 = (xor_ln896_42_fu_3829_p2 & tmp_139_reg_7293);

assign and_ln378_17_fu_4078_p2 = (xor_ln896_44_fu_4072_p2 & tmp_144_reg_7340);

assign and_ln378_18_fu_4321_p2 = (xor_ln896_46_fu_4315_p2 & tmp_149_reg_7387);

assign and_ln378_19_fu_4564_p2 = (xor_ln896_48_fu_4558_p2 & tmp_154_reg_7434);

assign and_ln378_1_fu_919_p2 = (xor_ln896_2_fu_913_p2 & tmp_79_reg_6729);

assign and_ln378_20_fu_4807_p2 = (xor_ln896_50_fu_4801_p2 & tmp_159_reg_7481);

assign and_ln378_21_fu_5050_p2 = (xor_ln896_52_fu_5044_p2 & tmp_164_reg_7528);

assign and_ln378_22_fu_5293_p2 = (xor_ln896_54_fu_5287_p2 & tmp_169_reg_7575);

assign and_ln378_23_fu_5536_p2 = (xor_ln896_56_fu_5530_p2 & tmp_174_reg_7622);

assign and_ln378_24_fu_5779_p2 = (xor_ln896_58_fu_5773_p2 & tmp_179_reg_7669);

assign and_ln378_25_fu_6009_p2 = (xor_ln896_60_fu_6003_p2 & tmp_184_reg_7716);

assign and_ln378_26_fu_6235_p2 = (xor_ln896_62_fu_6229_p2 & tmp_189_reg_7758);

assign and_ln378_3_fu_1162_p2 = (xor_ln896_5_fu_1156_p2 & tmp_84_reg_6776);

assign and_ln378_6_fu_1405_p2 = (xor_ln896_10_fu_1399_p2 & tmp_89_reg_6823);

assign and_ln378_7_fu_1648_p2 = (xor_ln896_16_fu_1642_p2 & tmp_94_reg_6870);

assign and_ln378_8_fu_1891_p2 = (xor_ln896_22_fu_1885_p2 & tmp_99_reg_6917);

assign and_ln378_9_fu_2134_p2 = (xor_ln896_27_fu_2128_p2 & tmp_104_reg_6964);

assign and_ln378_fu_676_p2 = (xor_ln896_fu_670_p2 & tmp_74_reg_6677);

assign and_ln890_10_fu_3147_p2 = (xor_ln890_16_fu_3141_p2 & icmp_ln1019_22_fu_3111_p2);

assign and_ln890_11_fu_3390_p2 = (xor_ln890_17_fu_3384_p2 & icmp_ln1019_24_fu_3354_p2);

assign and_ln890_12_fu_3633_p2 = (xor_ln890_18_fu_3627_p2 & icmp_ln1019_26_fu_3597_p2);

assign and_ln890_13_fu_3876_p2 = (xor_ln890_19_fu_3870_p2 & icmp_ln1019_28_fu_3840_p2);

assign and_ln890_14_fu_4119_p2 = (xor_ln890_20_fu_4113_p2 & icmp_ln1019_30_fu_4083_p2);

assign and_ln890_15_fu_4362_p2 = (xor_ln890_21_fu_4356_p2 & icmp_ln1019_32_fu_4326_p2);

assign and_ln890_16_fu_4605_p2 = (xor_ln890_22_fu_4599_p2 & icmp_ln1019_34_fu_4569_p2);

assign and_ln890_17_fu_4848_p2 = (xor_ln890_23_fu_4842_p2 & icmp_ln1019_36_fu_4812_p2);

assign and_ln890_18_fu_5091_p2 = (xor_ln890_24_fu_5085_p2 & icmp_ln1019_38_fu_5055_p2);

assign and_ln890_19_fu_5334_p2 = (xor_ln890_25_fu_5328_p2 & icmp_ln1019_40_fu_5298_p2);

assign and_ln890_1_fu_960_p2 = (xor_ln890_7_fu_954_p2 & icmp_ln1019_2_fu_924_p2);

assign and_ln890_20_fu_5577_p2 = (xor_ln890_26_fu_5571_p2 & icmp_ln1019_42_fu_5541_p2);

assign and_ln890_21_fu_5820_p2 = (xor_ln890_27_fu_5814_p2 & icmp_ln1019_44_fu_5784_p2);

assign and_ln890_22_fu_6050_p2 = (xor_ln890_28_fu_6044_p2 & icmp_ln1019_46_fu_6014_p2);

assign and_ln890_23_fu_6276_p2 = (xor_ln890_29_fu_6270_p2 & icmp_ln1019_48_fu_6240_p2);

assign and_ln890_2_fu_1203_p2 = (xor_ln890_8_fu_1197_p2 & icmp_ln1019_6_fu_1167_p2);

assign and_ln890_3_fu_1446_p2 = (xor_ln890_9_fu_1440_p2 & icmp_ln1019_8_fu_1410_p2);

assign and_ln890_4_fu_1689_p2 = (xor_ln890_10_fu_1683_p2 & icmp_ln1019_10_fu_1653_p2);

assign and_ln890_5_fu_1932_p2 = (xor_ln890_11_fu_1926_p2 & icmp_ln1019_12_fu_1896_p2);

assign and_ln890_6_fu_2175_p2 = (xor_ln890_12_fu_2169_p2 & icmp_ln1019_14_fu_2139_p2);

assign and_ln890_7_fu_2418_p2 = (xor_ln890_13_fu_2412_p2 & icmp_ln1019_16_fu_2382_p2);

assign and_ln890_8_fu_2661_p2 = (xor_ln890_14_fu_2655_p2 & icmp_ln1019_18_fu_2625_p2);

assign and_ln890_9_fu_2904_p2 = (xor_ln890_15_fu_2898_p2 & icmp_ln1019_20_fu_2868_p2);

assign and_ln890_fu_717_p2 = (xor_ln890_fu_711_p2 & icmp_ln1019_fu_681_p2);

assign and_ln891_10_fu_3161_p2 = (icmp_ln1019_23_fu_3116_p2 & and_ln378_13_fu_3106_p2);

assign and_ln891_11_fu_3404_p2 = (icmp_ln1019_25_fu_3359_p2 & and_ln378_14_fu_3349_p2);

assign and_ln891_12_fu_3647_p2 = (icmp_ln1019_27_fu_3602_p2 & and_ln378_15_fu_3592_p2);

assign and_ln891_13_fu_3890_p2 = (icmp_ln1019_29_fu_3845_p2 & and_ln378_16_fu_3835_p2);

assign and_ln891_14_fu_4133_p2 = (icmp_ln1019_31_fu_4088_p2 & and_ln378_17_fu_4078_p2);

assign and_ln891_15_fu_4376_p2 = (icmp_ln1019_33_fu_4331_p2 & and_ln378_18_fu_4321_p2);

assign and_ln891_16_fu_4619_p2 = (icmp_ln1019_35_fu_4574_p2 & and_ln378_19_fu_4564_p2);

assign and_ln891_17_fu_4862_p2 = (icmp_ln1019_37_fu_4817_p2 & and_ln378_20_fu_4807_p2);

assign and_ln891_18_fu_5105_p2 = (icmp_ln1019_39_fu_5060_p2 & and_ln378_21_fu_5050_p2);

assign and_ln891_19_fu_5348_p2 = (icmp_ln1019_41_fu_5303_p2 & and_ln378_22_fu_5293_p2);

assign and_ln891_1_fu_974_p2 = (icmp_ln1019_3_fu_929_p2 & and_ln378_1_fu_919_p2);

assign and_ln891_20_fu_5591_p2 = (icmp_ln1019_43_fu_5546_p2 & and_ln378_23_fu_5536_p2);

assign and_ln891_21_fu_5834_p2 = (icmp_ln1019_45_fu_5789_p2 & and_ln378_24_fu_5779_p2);

assign and_ln891_22_fu_6064_p2 = (icmp_ln1019_47_fu_6019_p2 & and_ln378_25_fu_6009_p2);

assign and_ln891_23_fu_6290_p2 = (icmp_ln1019_49_fu_6245_p2 & and_ln378_26_fu_6235_p2);

assign and_ln891_24_fu_1217_p2 = (icmp_ln1019_7_fu_1172_p2 & and_ln378_3_fu_1162_p2);

assign and_ln891_3_fu_1460_p2 = (icmp_ln1019_9_fu_1415_p2 & and_ln378_6_fu_1405_p2);

assign and_ln891_4_fu_1703_p2 = (icmp_ln1019_11_fu_1658_p2 & and_ln378_7_fu_1648_p2);

assign and_ln891_5_fu_1946_p2 = (icmp_ln1019_13_fu_1901_p2 & and_ln378_8_fu_1891_p2);

assign and_ln891_6_fu_2189_p2 = (icmp_ln1019_15_fu_2144_p2 & and_ln378_9_fu_2134_p2);

assign and_ln891_7_fu_2432_p2 = (icmp_ln1019_17_fu_2387_p2 & and_ln378_10_fu_2377_p2);

assign and_ln891_8_fu_2675_p2 = (icmp_ln1019_19_fu_2630_p2 & and_ln378_11_fu_2620_p2);

assign and_ln891_9_fu_2918_p2 = (icmp_ln1019_21_fu_2873_p2 & and_ln378_12_fu_2863_p2);

assign and_ln891_fu_731_p2 = (icmp_ln1019_1_fu_686_p2 & and_ln378_fu_676_p2);

assign and_ln895_10_fu_2455_p2 = (xor_ln895_22_fu_2450_p2 & or_ln895_7_fu_2444_p2);

assign and_ln895_11_fu_2698_p2 = (xor_ln895_24_fu_2693_p2 & or_ln895_8_fu_2687_p2);

assign and_ln895_12_fu_2941_p2 = (xor_ln895_26_fu_2936_p2 & or_ln895_9_fu_2930_p2);

assign and_ln895_13_fu_3184_p2 = (xor_ln895_28_fu_3179_p2 & or_ln895_10_fu_3173_p2);

assign and_ln895_14_fu_3427_p2 = (xor_ln895_30_fu_3422_p2 & or_ln895_11_fu_3416_p2);

assign and_ln895_15_fu_3670_p2 = (xor_ln895_32_fu_3665_p2 & or_ln895_12_fu_3659_p2);

assign and_ln895_16_fu_3913_p2 = (xor_ln895_34_fu_3908_p2 & or_ln895_13_fu_3902_p2);

assign and_ln895_17_fu_4156_p2 = (xor_ln895_36_fu_4151_p2 & or_ln895_14_fu_4145_p2);

assign and_ln895_18_fu_4399_p2 = (xor_ln895_38_fu_4394_p2 & or_ln895_15_fu_4388_p2);

assign and_ln895_19_fu_4642_p2 = (xor_ln895_40_fu_4637_p2 & or_ln895_16_fu_4631_p2);

assign and_ln895_1_fu_997_p2 = (xor_ln895_5_fu_992_p2 & or_ln895_1_fu_986_p2);

assign and_ln895_20_fu_4885_p2 = (xor_ln895_42_fu_4880_p2 & or_ln895_24_fu_4874_p2);

assign and_ln895_21_fu_5128_p2 = (xor_ln895_44_fu_5123_p2 & or_ln895_18_fu_5117_p2);

assign and_ln895_22_fu_5371_p2 = (xor_ln895_46_fu_5366_p2 & or_ln895_19_fu_5360_p2);

assign and_ln895_23_fu_5614_p2 = (xor_ln895_48_fu_5609_p2 & or_ln895_20_fu_5603_p2);

assign and_ln895_24_fu_5857_p2 = (xor_ln895_50_fu_5852_p2 & or_ln895_21_fu_5846_p2);

assign and_ln895_25_fu_6087_p2 = (xor_ln895_52_fu_6082_p2 & or_ln895_22_fu_6076_p2);

assign and_ln895_26_fu_6313_p2 = (xor_ln895_54_fu_6308_p2 & or_ln895_23_fu_6302_p2);

assign and_ln895_3_fu_1240_p2 = (xor_ln895_11_fu_1235_p2 & or_ln895_17_fu_1229_p2);

assign and_ln895_6_fu_1483_p2 = (xor_ln895_14_fu_1478_p2 & or_ln895_3_fu_1472_p2);

assign and_ln895_7_fu_1726_p2 = (xor_ln895_16_fu_1721_p2 & or_ln895_4_fu_1715_p2);

assign and_ln895_8_fu_1969_p2 = (xor_ln895_18_fu_1964_p2 & or_ln895_5_fu_1958_p2);

assign and_ln895_9_fu_2212_p2 = (xor_ln895_20_fu_2207_p2 & or_ln895_6_fu_2201_p2);

assign and_ln895_fu_754_p2 = (xor_ln895_3_fu_749_p2 & or_ln895_fu_743_p2);

assign and_ln896_10_fu_2479_p2 = (xor_ln896_66_fu_2473_p2 & tmp_108_reg_7000);

assign and_ln896_11_fu_2722_p2 = (xor_ln896_67_fu_2716_p2 & tmp_113_reg_7047);

assign and_ln896_12_fu_2965_p2 = (xor_ln896_68_fu_2959_p2 & tmp_118_reg_7094);

assign and_ln896_13_fu_3208_p2 = (xor_ln896_69_fu_3202_p2 & tmp_123_reg_7141);

assign and_ln896_14_fu_3451_p2 = (xor_ln896_70_fu_3445_p2 & tmp_128_reg_7188);

assign and_ln896_15_fu_3694_p2 = (xor_ln896_71_fu_3688_p2 & tmp_133_reg_7235);

assign and_ln896_16_fu_3937_p2 = (xor_ln896_72_fu_3931_p2 & tmp_138_reg_7282);

assign and_ln896_17_fu_4180_p2 = (xor_ln896_73_fu_4174_p2 & tmp_143_reg_7329);

assign and_ln896_18_fu_4423_p2 = (xor_ln896_74_fu_4417_p2 & tmp_148_reg_7376);

assign and_ln896_19_fu_4666_p2 = (xor_ln896_75_fu_4660_p2 & tmp_153_reg_7423);

assign and_ln896_1_fu_1021_p2 = (xor_ln896_23_fu_1015_p2 & tmp_78_reg_6718);

assign and_ln896_20_fu_4909_p2 = (xor_ln896_76_fu_4903_p2 & tmp_158_reg_7470);

assign and_ln896_21_fu_5152_p2 = (xor_ln896_77_fu_5146_p2 & tmp_163_reg_7517);

assign and_ln896_22_fu_5395_p2 = (xor_ln896_78_fu_5389_p2 & tmp_168_reg_7564);

assign and_ln896_23_fu_5638_p2 = (xor_ln896_79_fu_5632_p2 & tmp_173_reg_7611);

assign and_ln896_24_fu_5881_p2 = (xor_ln896_80_fu_5875_p2 & tmp_178_reg_7658);

assign and_ln896_25_fu_6111_p2 = (xor_ln896_81_fu_6105_p2 & tmp_183_reg_7705);

assign and_ln896_26_fu_6337_p2 = (xor_ln896_82_fu_6331_p2 & tmp_188_reg_7747);

assign and_ln896_3_fu_1264_p2 = (xor_ln896_24_fu_1258_p2 & tmp_83_reg_6765);

assign and_ln896_6_fu_1507_p2 = (xor_ln896_25_fu_1501_p2 & tmp_88_reg_6812);

assign and_ln896_7_fu_1750_p2 = (xor_ln896_28_fu_1744_p2 & tmp_93_reg_6859);

assign and_ln896_8_fu_1993_p2 = (xor_ln896_64_fu_1987_p2 & tmp_98_reg_6906);

assign and_ln896_9_fu_2236_p2 = (xor_ln896_65_fu_2230_p2 & tmp_103_reg_6953);

assign and_ln896_fu_778_p2 = (xor_ln896_20_fu_772_p2 & tmp_73_reg_6666);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage0_iter24 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage0_iter25 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

assign icmp_ln1019_10_fu_1653_p2 = ((tmp_12_reg_6875 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_11_fu_1658_p2 = ((tmp_13_reg_6880 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_12_fu_1896_p2 = ((tmp_15_reg_6922 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_13_fu_1901_p2 = ((tmp_16_reg_6927 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_14_fu_2139_p2 = ((tmp_18_reg_6969 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_15_fu_2144_p2 = ((tmp_19_reg_6974 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_16_fu_2382_p2 = ((tmp_21_reg_7016 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_17_fu_2387_p2 = ((tmp_22_reg_7021 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_18_fu_2625_p2 = ((tmp_24_reg_7063 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_19_fu_2630_p2 = ((tmp_25_reg_7068 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_1_fu_686_p2 = ((tmp_2_reg_6692 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_20_fu_2868_p2 = ((tmp_27_reg_7110 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_21_fu_2873_p2 = ((tmp_28_reg_7115 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_22_fu_3111_p2 = ((tmp_30_reg_7157 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_23_fu_3116_p2 = ((tmp_31_reg_7162 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_24_fu_3354_p2 = ((tmp_33_reg_7204 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_25_fu_3359_p2 = ((tmp_34_reg_7209 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_26_fu_3597_p2 = ((tmp_36_reg_7251 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_27_fu_3602_p2 = ((tmp_37_reg_7256 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_28_fu_3840_p2 = ((tmp_39_reg_7298 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_29_fu_3845_p2 = ((tmp_40_reg_7303 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_2_fu_924_p2 = ((tmp_4_reg_6734 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_30_fu_4083_p2 = ((tmp_42_reg_7345 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_31_fu_4088_p2 = ((tmp_43_reg_7350 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_32_fu_4326_p2 = ((tmp_45_reg_7392 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_33_fu_4331_p2 = ((tmp_46_reg_7397 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_34_fu_4569_p2 = ((tmp_48_reg_7439 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_35_fu_4574_p2 = ((tmp_49_reg_7444 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_36_fu_4812_p2 = ((tmp_51_reg_7486 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_37_fu_4817_p2 = ((tmp_52_reg_7491 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_38_fu_5055_p2 = ((tmp_54_reg_7533 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_39_fu_5060_p2 = ((tmp_55_reg_7538 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_3_fu_929_p2 = ((tmp_5_reg_6739 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_40_fu_5298_p2 = ((tmp_57_reg_7580 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_41_fu_5303_p2 = ((tmp_58_reg_7585 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_42_fu_5541_p2 = ((tmp_60_reg_7627 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_43_fu_5546_p2 = ((tmp_61_reg_7632 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_44_fu_5784_p2 = ((tmp_63_reg_7674 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_45_fu_5789_p2 = ((tmp_64_reg_7679 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_46_fu_6014_p2 = ((tmp_66_reg_7721 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_47_fu_6019_p2 = ((tmp_67_reg_7726 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_48_fu_6240_p2 = ((tmp_69_reg_7763 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_49_fu_6245_p2 = ((tmp_70_reg_7768 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_6_fu_1167_p2 = ((tmp_7_reg_6781 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_7_fu_1172_p2 = ((tmp_8_reg_6786 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_8_fu_1410_p2 = ((tmp_10_reg_6828 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1019_9_fu_1415_p2 = ((tmp_11_reg_6833 == 16'd65535) ? 1'b1 : 1'b0);

assign icmp_ln1019_fu_681_p2 = ((tmp_1_reg_6687 == 15'd32767) ? 1'b1 : 1'b0);

assign icmp_ln1420_1_fu_6369_p2 = ((trunc_ln25_reg_6622_pp0_iter24_reg == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln1420_2_fu_6374_p2 = ((trunc_ln25_reg_6622_pp0_iter24_reg == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln1420_fu_6364_p2 = ((trunc_ln25_reg_6622_pp0_iter24_reg == 2'd0) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_514_p2 = ((ap_sig_allocacmp_i == 3'd4) ? 1'b1 : 1'b0);

assign icmp_ln878_10_fu_2878_p2 = ((tmp_28_reg_7115 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_11_fu_3121_p2 = ((tmp_31_reg_7162 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_12_fu_3364_p2 = ((tmp_34_reg_7209 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_13_fu_3607_p2 = ((tmp_37_reg_7256 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_14_fu_3850_p2 = ((tmp_40_reg_7303 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_15_fu_4093_p2 = ((tmp_43_reg_7350 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_16_fu_4336_p2 = ((tmp_46_reg_7397 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_17_fu_4579_p2 = ((tmp_49_reg_7444 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_18_fu_4822_p2 = ((tmp_52_reg_7491 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_19_fu_5065_p2 = ((tmp_55_reg_7538 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_1_fu_934_p2 = ((tmp_5_reg_6739 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_20_fu_5308_p2 = ((tmp_58_reg_7585 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_21_fu_5551_p2 = ((tmp_61_reg_7632 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_22_fu_5794_p2 = ((tmp_64_reg_7679 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_23_fu_6024_p2 = ((tmp_67_reg_7726 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_24_fu_6250_p2 = ((tmp_70_reg_7768 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_3_fu_1177_p2 = ((tmp_8_reg_6786 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_4_fu_1420_p2 = ((tmp_11_reg_6833 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_5_fu_1663_p2 = ((tmp_13_reg_6880 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_6_fu_1906_p2 = ((tmp_16_reg_6927 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_7_fu_2149_p2 = ((tmp_19_reg_6974 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_8_fu_2392_p2 = ((tmp_22_reg_7021 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_9_fu_2635_p2 = ((tmp_25_reg_7068 == 16'd0) ? 1'b1 : 1'b0);

assign icmp_ln878_fu_691_p2 = ((tmp_2_reg_6692 == 16'd0) ? 1'b1 : 1'b0);

assign mul_ln1273_10_fu_2086_p0 = sext_ln1273_7_cast_reg_6578;

assign mul_ln1273_11_fu_2329_p0 = sext_ln1273_8_cast_reg_6573;

assign mul_ln1273_12_fu_2572_p0 = sext_ln1273_9_cast_reg_6568;

assign mul_ln1273_13_fu_2815_p0 = sext_ln1273_10_cast_reg_6563;

assign mul_ln1273_14_fu_3058_p0 = sext_ln1273_11_cast_reg_6558;

assign mul_ln1273_15_fu_3301_p0 = sext_ln1273_12_cast_reg_6553;

assign mul_ln1273_16_fu_3544_p0 = sext_ln1273_13_cast_reg_6548;

assign mul_ln1273_17_fu_3787_p0 = sext_ln1273_14_cast_reg_6543;

assign mul_ln1273_18_fu_4030_p0 = sext_ln1273_15_cast_reg_6538;

assign mul_ln1273_19_fu_4273_p0 = sext_ln1273_16_cast_reg_6533;

assign mul_ln1273_1_fu_628_p0 = sext_ln1273_1_cast_reg_6608;

assign mul_ln1273_20_fu_4516_p0 = sext_ln1273_17_cast_reg_6528;

assign mul_ln1273_21_fu_4759_p0 = sext_ln1273_18_cast_reg_6523;

assign mul_ln1273_22_fu_5002_p0 = sext_ln1273_19_cast_reg_6518;

assign mul_ln1273_23_fu_5245_p0 = sext_ln1273_20_cast_reg_6513;

assign mul_ln1273_24_fu_5488_p0 = sext_ln1273_21_cast_reg_6508;

assign mul_ln1273_25_fu_5731_p0 = sext_ln1273_22_cast_reg_6503;

assign mul_ln1273_26_fu_5974_p0 = sext_ln1273_23_cast_reg_6498;

assign mul_ln1273_3_fu_871_p0 = sext_ln1273_24_cast_reg_6603;

assign mul_ln1273_6_fu_1114_p0 = sext_ln1273_3_cast_reg_6598;

assign mul_ln1273_7_fu_1357_p0 = sext_ln1273_4_cast_reg_6593;

assign mul_ln1273_8_fu_1600_p0 = sext_ln1273_5_cast_reg_6588;

assign mul_ln1273_9_fu_1843_p0 = sext_ln1273_6_cast_reg_6583;

assign mul_ln1273_fu_566_p0 = sext_ln1273_cast_reg_6613;

assign or_ln1420_1_fu_6385_p2 = (or_ln1420_fu_6379_p2 | icmp_ln1420_fu_6364_p2);

assign or_ln1420_fu_6379_p2 = (icmp_ln1420_2_fu_6374_p2 | icmp_ln1420_1_fu_6369_p2);

assign or_ln346_10_fu_2484_p2 = (and_ln896_10_fu_2479_p2 | and_ln895_10_fu_2455_p2);

assign or_ln346_11_fu_2727_p2 = (and_ln896_11_fu_2722_p2 | and_ln895_11_fu_2698_p2);

assign or_ln346_12_fu_2970_p2 = (and_ln896_12_fu_2965_p2 | and_ln895_12_fu_2941_p2);

assign or_ln346_13_fu_3213_p2 = (and_ln896_13_fu_3208_p2 | and_ln895_13_fu_3184_p2);

assign or_ln346_14_fu_3456_p2 = (and_ln896_14_fu_3451_p2 | and_ln895_14_fu_3427_p2);

assign or_ln346_15_fu_3699_p2 = (and_ln896_15_fu_3694_p2 | and_ln895_15_fu_3670_p2);

assign or_ln346_16_fu_3942_p2 = (and_ln896_16_fu_3937_p2 | and_ln895_16_fu_3913_p2);

assign or_ln346_17_fu_4185_p2 = (and_ln896_17_fu_4180_p2 | and_ln895_17_fu_4156_p2);

assign or_ln346_18_fu_4428_p2 = (and_ln896_18_fu_4423_p2 | and_ln895_18_fu_4399_p2);

assign or_ln346_19_fu_4671_p2 = (and_ln896_19_fu_4666_p2 | and_ln895_19_fu_4642_p2);

assign or_ln346_1_fu_1026_p2 = (and_ln896_1_fu_1021_p2 | and_ln895_1_fu_997_p2);

assign or_ln346_20_fu_4914_p2 = (and_ln896_20_fu_4909_p2 | and_ln895_20_fu_4885_p2);

assign or_ln346_21_fu_5157_p2 = (and_ln896_21_fu_5152_p2 | and_ln895_21_fu_5128_p2);

assign or_ln346_22_fu_5400_p2 = (and_ln896_22_fu_5395_p2 | and_ln895_22_fu_5371_p2);

assign or_ln346_23_fu_5643_p2 = (and_ln896_23_fu_5638_p2 | and_ln895_23_fu_5614_p2);

assign or_ln346_24_fu_5886_p2 = (and_ln896_24_fu_5881_p2 | and_ln895_24_fu_5857_p2);

assign or_ln346_25_fu_6116_p2 = (and_ln896_25_fu_6111_p2 | and_ln895_25_fu_6087_p2);

assign or_ln346_26_fu_6350_p2 = (and_ln896_26_fu_6337_p2 | and_ln895_26_fu_6313_p2);

assign or_ln346_3_fu_1269_p2 = (and_ln896_3_fu_1264_p2 | and_ln895_3_fu_1240_p2);

assign or_ln346_6_fu_1512_p2 = (and_ln896_6_fu_1507_p2 | and_ln895_6_fu_1483_p2);

assign or_ln346_7_fu_1755_p2 = (and_ln896_7_fu_1750_p2 | and_ln895_7_fu_1726_p2);

assign or_ln346_8_fu_1998_p2 = (and_ln896_8_fu_1993_p2 | and_ln895_8_fu_1969_p2);

assign or_ln346_9_fu_2241_p2 = (and_ln896_9_fu_2236_p2 | and_ln895_9_fu_2212_p2);

assign or_ln346_fu_783_p2 = (and_ln896_fu_778_p2 | and_ln895_fu_754_p2);

assign or_ln895_10_fu_3173_p2 = (xor_ln895_27_fu_3167_p2 | tmp_126_fu_3092_p3);

assign or_ln895_11_fu_3416_p2 = (xor_ln895_29_fu_3410_p2 | tmp_131_fu_3335_p3);

assign or_ln895_12_fu_3659_p2 = (xor_ln895_31_fu_3653_p2 | tmp_136_fu_3578_p3);

assign or_ln895_13_fu_3902_p2 = (xor_ln895_33_fu_3896_p2 | tmp_141_fu_3821_p3);

assign or_ln895_14_fu_4145_p2 = (xor_ln895_35_fu_4139_p2 | tmp_146_fu_4064_p3);

assign or_ln895_15_fu_4388_p2 = (xor_ln895_37_fu_4382_p2 | tmp_151_fu_4307_p3);

assign or_ln895_16_fu_4631_p2 = (xor_ln895_39_fu_4625_p2 | tmp_156_fu_4550_p3);

assign or_ln895_17_fu_1229_p2 = (xor_ln895_10_fu_1223_p2 | tmp_86_fu_1148_p3);

assign or_ln895_18_fu_5117_p2 = (xor_ln895_43_fu_5111_p2 | tmp_166_fu_5036_p3);

assign or_ln895_19_fu_5360_p2 = (xor_ln895_45_fu_5354_p2 | tmp_171_fu_5279_p3);

assign or_ln895_1_fu_986_p2 = (xor_ln895_4_fu_980_p2 | tmp_81_fu_905_p3);

assign or_ln895_20_fu_5603_p2 = (xor_ln895_47_fu_5597_p2 | tmp_176_fu_5522_p3);

assign or_ln895_21_fu_5846_p2 = (xor_ln895_49_fu_5840_p2 | tmp_181_fu_5765_p3);

assign or_ln895_22_fu_6076_p2 = (xor_ln895_51_fu_6070_p2 | tmp_186_fu_5995_p3);

assign or_ln895_23_fu_6302_p2 = (xor_ln895_53_fu_6296_p2 | tmp_191_fu_6221_p3);

assign or_ln895_24_fu_4874_p2 = (xor_ln895_41_fu_4868_p2 | tmp_161_fu_4793_p3);

assign or_ln895_3_fu_1472_p2 = (xor_ln895_fu_1466_p2 | tmp_91_fu_1391_p3);

assign or_ln895_4_fu_1715_p2 = (xor_ln895_15_fu_1709_p2 | tmp_96_fu_1634_p3);

assign or_ln895_5_fu_1958_p2 = (xor_ln895_17_fu_1952_p2 | tmp_101_fu_1877_p3);

assign or_ln895_6_fu_2201_p2 = (xor_ln895_19_fu_2195_p2 | tmp_106_fu_2120_p3);

assign or_ln895_7_fu_2444_p2 = (xor_ln895_21_fu_2438_p2 | tmp_111_fu_2363_p3);

assign or_ln895_8_fu_2687_p2 = (xor_ln895_23_fu_2681_p2 | tmp_116_fu_2606_p3);

assign or_ln895_9_fu_2930_p2 = (xor_ln895_25_fu_2924_p2 | tmp_121_fu_2849_p3);

assign or_ln895_fu_743_p2 = (xor_ln895_2_fu_737_p2 | tmp_76_fu_662_p3);

assign or_ln896_10_fu_3196_p2 = (xor_ln896_37_fu_3190_p2 | xor_ln896_36_fu_3100_p2);

assign or_ln896_11_fu_3439_p2 = (xor_ln896_39_fu_3433_p2 | xor_ln896_38_fu_3343_p2);

assign or_ln896_12_fu_3682_p2 = (xor_ln896_41_fu_3676_p2 | xor_ln896_40_fu_3586_p2);

assign or_ln896_13_fu_3925_p2 = (xor_ln896_43_fu_3919_p2 | xor_ln896_42_fu_3829_p2);

assign or_ln896_14_fu_4168_p2 = (xor_ln896_45_fu_4162_p2 | xor_ln896_44_fu_4072_p2);

assign or_ln896_15_fu_4411_p2 = (xor_ln896_47_fu_4405_p2 | xor_ln896_46_fu_4315_p2);

assign or_ln896_16_fu_4654_p2 = (xor_ln896_49_fu_4648_p2 | xor_ln896_48_fu_4558_p2);

assign or_ln896_17_fu_4897_p2 = (xor_ln896_51_fu_4891_p2 | xor_ln896_50_fu_4801_p2);

assign or_ln896_18_fu_1252_p2 = (xor_ln896_9_fu_1246_p2 | xor_ln896_5_fu_1156_p2);

assign or_ln896_19_fu_5383_p2 = (xor_ln896_55_fu_5377_p2 | xor_ln896_54_fu_5287_p2);

assign or_ln896_1_fu_1009_p2 = (xor_ln896_4_fu_1003_p2 | xor_ln896_2_fu_913_p2);

assign or_ln896_20_fu_5626_p2 = (xor_ln896_57_fu_5620_p2 | xor_ln896_56_fu_5530_p2);

assign or_ln896_21_fu_5869_p2 = (xor_ln896_59_fu_5863_p2 | xor_ln896_58_fu_5773_p2);

assign or_ln896_22_fu_6099_p2 = (xor_ln896_61_fu_6093_p2 | xor_ln896_60_fu_6003_p2);

assign or_ln896_23_fu_6325_p2 = (xor_ln896_63_fu_6319_p2 | xor_ln896_62_fu_6229_p2);

assign or_ln896_24_fu_5140_p2 = (xor_ln896_53_fu_5134_p2 | xor_ln896_52_fu_5044_p2);

assign or_ln896_3_fu_1495_p2 = (xor_ln896_15_fu_1489_p2 | xor_ln896_10_fu_1399_p2);

assign or_ln896_4_fu_1738_p2 = (xor_ln896_21_fu_1732_p2 | xor_ln896_16_fu_1642_p2);

assign or_ln896_5_fu_1981_p2 = (xor_ln896_26_fu_1975_p2 | xor_ln896_22_fu_1885_p2);

assign or_ln896_6_fu_2224_p2 = (xor_ln896_29_fu_2218_p2 | xor_ln896_27_fu_2128_p2);

assign or_ln896_7_fu_2467_p2 = (xor_ln896_31_fu_2461_p2 | xor_ln896_30_fu_2371_p2);

assign or_ln896_8_fu_2710_p2 = (xor_ln896_33_fu_2704_p2 | xor_ln896_32_fu_2614_p2);

assign or_ln896_9_fu_2953_p2 = (xor_ln896_35_fu_2947_p2 | xor_ln896_34_fu_2857_p2);

assign or_ln896_fu_766_p2 = (xor_ln896_fu_670_p2 | xor_ln896_1_fu_760_p2);

assign select_ln346_10_fu_1761_p3 = ((and_ln895_7_fu_1726_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_11_fu_1769_p3 = ((or_ln346_7_fu_1755_p2[0:0] == 1'b1) ? select_ln346_10_fu_1761_p3 : add_ln377_7_fu_1629_p2);

assign select_ln346_12_fu_2004_p3 = ((and_ln895_8_fu_1969_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_13_fu_2012_p3 = ((or_ln346_8_fu_1998_p2[0:0] == 1'b1) ? select_ln346_12_fu_2004_p3 : add_ln377_8_fu_1872_p2);

assign select_ln346_14_fu_2247_p3 = ((and_ln895_9_fu_2212_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_15_fu_2490_p3 = ((and_ln895_10_fu_2455_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_16_fu_2498_p3 = ((or_ln346_10_fu_2484_p2[0:0] == 1'b1) ? select_ln346_15_fu_2490_p3 : add_ln377_10_fu_2358_p2);

assign select_ln346_17_fu_2733_p3 = ((and_ln895_11_fu_2698_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_18_fu_2741_p3 = ((or_ln346_11_fu_2727_p2[0:0] == 1'b1) ? select_ln346_17_fu_2733_p3 : add_ln377_11_fu_2601_p2);

assign select_ln346_19_fu_2976_p3 = ((and_ln895_12_fu_2941_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_20_fu_2984_p3 = ((or_ln346_12_fu_2970_p2[0:0] == 1'b1) ? select_ln346_19_fu_2976_p3 : add_ln377_12_fu_2844_p2);

assign select_ln346_21_fu_3219_p3 = ((and_ln895_13_fu_3184_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_22_fu_3227_p3 = ((or_ln346_13_fu_3213_p2[0:0] == 1'b1) ? select_ln346_21_fu_3219_p3 : add_ln377_13_fu_3087_p2);

assign select_ln346_23_fu_3462_p3 = ((and_ln895_14_fu_3427_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_24_fu_3470_p3 = ((or_ln346_14_fu_3456_p2[0:0] == 1'b1) ? select_ln346_23_fu_3462_p3 : add_ln377_14_fu_3330_p2);

assign select_ln346_25_fu_3705_p3 = ((and_ln895_15_fu_3670_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_26_fu_3713_p3 = ((or_ln346_15_fu_3699_p2[0:0] == 1'b1) ? select_ln346_25_fu_3705_p3 : add_ln377_15_fu_3573_p2);

assign select_ln346_27_fu_3948_p3 = ((and_ln895_16_fu_3913_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_28_fu_3956_p3 = ((or_ln346_16_fu_3942_p2[0:0] == 1'b1) ? select_ln346_27_fu_3948_p3 : add_ln377_16_fu_3816_p2);

assign select_ln346_29_fu_4191_p3 = ((and_ln895_17_fu_4156_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_2_fu_789_p3 = ((and_ln895_fu_754_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_30_fu_4199_p3 = ((or_ln346_17_fu_4185_p2[0:0] == 1'b1) ? select_ln346_29_fu_4191_p3 : add_ln377_17_fu_4059_p2);

assign select_ln346_31_fu_4434_p3 = ((and_ln895_18_fu_4399_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_32_fu_4442_p3 = ((or_ln346_18_fu_4428_p2[0:0] == 1'b1) ? select_ln346_31_fu_4434_p3 : add_ln377_18_fu_4302_p2);

assign select_ln346_33_fu_4677_p3 = ((and_ln895_19_fu_4642_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_34_fu_4685_p3 = ((or_ln346_19_fu_4671_p2[0:0] == 1'b1) ? select_ln346_33_fu_4677_p3 : add_ln377_19_fu_4545_p2);

assign select_ln346_35_fu_4920_p3 = ((and_ln895_20_fu_4885_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_36_fu_4928_p3 = ((or_ln346_20_fu_4914_p2[0:0] == 1'b1) ? select_ln346_35_fu_4920_p3 : add_ln377_20_fu_4788_p2);

assign select_ln346_37_fu_5163_p3 = ((and_ln895_21_fu_5128_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_38_fu_5171_p3 = ((or_ln346_21_fu_5157_p2[0:0] == 1'b1) ? select_ln346_37_fu_5163_p3 : add_ln377_21_fu_5031_p2);

assign select_ln346_39_fu_5406_p3 = ((and_ln895_22_fu_5371_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_3_fu_797_p3 = ((or_ln346_fu_783_p2[0:0] == 1'b1) ? select_ln346_2_fu_789_p3 : add_ln377_fu_657_p2);

assign select_ln346_40_fu_5414_p3 = ((or_ln346_22_fu_5400_p2[0:0] == 1'b1) ? select_ln346_39_fu_5406_p3 : add_ln377_22_fu_5274_p2);

assign select_ln346_41_fu_5649_p3 = ((and_ln895_23_fu_5614_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_42_fu_5657_p3 = ((or_ln346_23_fu_5643_p2[0:0] == 1'b1) ? select_ln346_41_fu_5649_p3 : add_ln377_23_fu_5517_p2);

assign select_ln346_43_fu_5892_p3 = ((and_ln895_24_fu_5857_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_44_fu_5900_p3 = ((or_ln346_24_fu_5886_p2[0:0] == 1'b1) ? select_ln346_43_fu_5892_p3 : add_ln377_24_fu_5760_p2);

assign select_ln346_45_fu_6122_p3 = ((and_ln895_25_fu_6087_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_46_fu_6130_p3 = ((or_ln346_25_fu_6116_p2[0:0] == 1'b1) ? select_ln346_45_fu_6122_p3 : add_ln377_25_fu_5990_p2);

assign select_ln346_47_fu_6342_p3 = ((and_ln895_26_fu_6313_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_4_fu_1032_p3 = ((and_ln895_1_fu_997_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_5_fu_1040_p3 = ((or_ln346_1_fu_1026_p2[0:0] == 1'b1) ? select_ln346_4_fu_1032_p3 : add_ln377_1_fu_900_p2);

assign select_ln346_6_fu_1275_p3 = ((and_ln895_3_fu_1240_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_7_fu_1283_p3 = ((or_ln346_3_fu_1269_p2[0:0] == 1'b1) ? select_ln346_6_fu_1275_p3 : add_ln377_3_fu_1143_p2);

assign select_ln346_8_fu_1518_p3 = ((and_ln895_6_fu_1483_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_9_fu_1526_p3 = ((or_ln346_6_fu_1512_p2[0:0] == 1'b1) ? select_ln346_8_fu_1518_p3 : add_ln377_6_fu_1386_p2);

assign select_ln346_fu_2255_p3 = ((or_ln346_9_fu_2241_p2[0:0] == 1'b1) ? select_ln346_14_fu_2247_p3 : add_ln377_9_fu_2115_p2);

assign select_ln888_10_fu_2883_p3 = ((and_ln378_12_fu_2863_p2[0:0] == 1'b1) ? icmp_ln1019_21_fu_2873_p2 : icmp_ln878_10_fu_2878_p2);

assign select_ln888_11_fu_3126_p3 = ((and_ln378_13_fu_3106_p2[0:0] == 1'b1) ? icmp_ln1019_23_fu_3116_p2 : icmp_ln878_11_fu_3121_p2);

assign select_ln888_12_fu_3369_p3 = ((and_ln378_14_fu_3349_p2[0:0] == 1'b1) ? icmp_ln1019_25_fu_3359_p2 : icmp_ln878_12_fu_3364_p2);

assign select_ln888_13_fu_3612_p3 = ((and_ln378_15_fu_3592_p2[0:0] == 1'b1) ? icmp_ln1019_27_fu_3602_p2 : icmp_ln878_13_fu_3607_p2);

assign select_ln888_14_fu_3855_p3 = ((and_ln378_16_fu_3835_p2[0:0] == 1'b1) ? icmp_ln1019_29_fu_3845_p2 : icmp_ln878_14_fu_3850_p2);

assign select_ln888_15_fu_4098_p3 = ((and_ln378_17_fu_4078_p2[0:0] == 1'b1) ? icmp_ln1019_31_fu_4088_p2 : icmp_ln878_15_fu_4093_p2);

assign select_ln888_16_fu_4341_p3 = ((and_ln378_18_fu_4321_p2[0:0] == 1'b1) ? icmp_ln1019_33_fu_4331_p2 : icmp_ln878_16_fu_4336_p2);

assign select_ln888_17_fu_4584_p3 = ((and_ln378_19_fu_4564_p2[0:0] == 1'b1) ? icmp_ln1019_35_fu_4574_p2 : icmp_ln878_17_fu_4579_p2);

assign select_ln888_18_fu_4827_p3 = ((and_ln378_20_fu_4807_p2[0:0] == 1'b1) ? icmp_ln1019_37_fu_4817_p2 : icmp_ln878_18_fu_4822_p2);

assign select_ln888_19_fu_5070_p3 = ((and_ln378_21_fu_5050_p2[0:0] == 1'b1) ? icmp_ln1019_39_fu_5060_p2 : icmp_ln878_19_fu_5065_p2);

assign select_ln888_1_fu_939_p3 = ((and_ln378_1_fu_919_p2[0:0] == 1'b1) ? icmp_ln1019_3_fu_929_p2 : icmp_ln878_1_fu_934_p2);

assign select_ln888_20_fu_5313_p3 = ((and_ln378_22_fu_5293_p2[0:0] == 1'b1) ? icmp_ln1019_41_fu_5303_p2 : icmp_ln878_20_fu_5308_p2);

assign select_ln888_21_fu_5556_p3 = ((and_ln378_23_fu_5536_p2[0:0] == 1'b1) ? icmp_ln1019_43_fu_5546_p2 : icmp_ln878_21_fu_5551_p2);

assign select_ln888_22_fu_5799_p3 = ((and_ln378_24_fu_5779_p2[0:0] == 1'b1) ? icmp_ln1019_45_fu_5789_p2 : icmp_ln878_22_fu_5794_p2);

assign select_ln888_23_fu_6029_p3 = ((and_ln378_25_fu_6009_p2[0:0] == 1'b1) ? icmp_ln1019_47_fu_6019_p2 : icmp_ln878_23_fu_6024_p2);

assign select_ln888_24_fu_6255_p3 = ((and_ln378_26_fu_6235_p2[0:0] == 1'b1) ? icmp_ln1019_49_fu_6245_p2 : icmp_ln878_24_fu_6250_p2);

assign select_ln888_3_fu_1182_p3 = ((and_ln378_3_fu_1162_p2[0:0] == 1'b1) ? icmp_ln1019_7_fu_1172_p2 : icmp_ln878_3_fu_1177_p2);

assign select_ln888_4_fu_1425_p3 = ((and_ln378_6_fu_1405_p2[0:0] == 1'b1) ? icmp_ln1019_9_fu_1415_p2 : icmp_ln878_4_fu_1420_p2);

assign select_ln888_5_fu_1668_p3 = ((and_ln378_7_fu_1648_p2[0:0] == 1'b1) ? icmp_ln1019_11_fu_1658_p2 : icmp_ln878_5_fu_1663_p2);

assign select_ln888_6_fu_1911_p3 = ((and_ln378_8_fu_1891_p2[0:0] == 1'b1) ? icmp_ln1019_13_fu_1901_p2 : icmp_ln878_6_fu_1906_p2);

assign select_ln888_7_fu_2154_p3 = ((and_ln378_9_fu_2134_p2[0:0] == 1'b1) ? icmp_ln1019_15_fu_2144_p2 : icmp_ln878_7_fu_2149_p2);

assign select_ln888_8_fu_2397_p3 = ((and_ln378_10_fu_2377_p2[0:0] == 1'b1) ? icmp_ln1019_17_fu_2387_p2 : icmp_ln878_8_fu_2392_p2);

assign select_ln888_9_fu_2640_p3 = ((and_ln378_11_fu_2620_p2[0:0] == 1'b1) ? icmp_ln1019_19_fu_2630_p2 : icmp_ln878_9_fu_2635_p2);

assign select_ln888_fu_696_p3 = ((and_ln378_fu_676_p2[0:0] == 1'b1) ? icmp_ln1019_1_fu_686_p2 : icmp_ln878_fu_691_p2);

assign select_ln890_10_fu_2910_p3 = ((and_ln378_12_fu_2863_p2[0:0] == 1'b1) ? and_ln890_9_fu_2904_p2 : icmp_ln1019_21_fu_2873_p2);

assign select_ln890_11_fu_3153_p3 = ((and_ln378_13_fu_3106_p2[0:0] == 1'b1) ? and_ln890_10_fu_3147_p2 : icmp_ln1019_23_fu_3116_p2);

assign select_ln890_12_fu_3396_p3 = ((and_ln378_14_fu_3349_p2[0:0] == 1'b1) ? and_ln890_11_fu_3390_p2 : icmp_ln1019_25_fu_3359_p2);

assign select_ln890_13_fu_3639_p3 = ((and_ln378_15_fu_3592_p2[0:0] == 1'b1) ? and_ln890_12_fu_3633_p2 : icmp_ln1019_27_fu_3602_p2);

assign select_ln890_14_fu_3882_p3 = ((and_ln378_16_fu_3835_p2[0:0] == 1'b1) ? and_ln890_13_fu_3876_p2 : icmp_ln1019_29_fu_3845_p2);

assign select_ln890_15_fu_4125_p3 = ((and_ln378_17_fu_4078_p2[0:0] == 1'b1) ? and_ln890_14_fu_4119_p2 : icmp_ln1019_31_fu_4088_p2);

assign select_ln890_16_fu_4368_p3 = ((and_ln378_18_fu_4321_p2[0:0] == 1'b1) ? and_ln890_15_fu_4362_p2 : icmp_ln1019_33_fu_4331_p2);

assign select_ln890_17_fu_4611_p3 = ((and_ln378_19_fu_4564_p2[0:0] == 1'b1) ? and_ln890_16_fu_4605_p2 : icmp_ln1019_35_fu_4574_p2);

assign select_ln890_18_fu_4854_p3 = ((and_ln378_20_fu_4807_p2[0:0] == 1'b1) ? and_ln890_17_fu_4848_p2 : icmp_ln1019_37_fu_4817_p2);

assign select_ln890_19_fu_5097_p3 = ((and_ln378_21_fu_5050_p2[0:0] == 1'b1) ? and_ln890_18_fu_5091_p2 : icmp_ln1019_39_fu_5060_p2);

assign select_ln890_1_fu_966_p3 = ((and_ln378_1_fu_919_p2[0:0] == 1'b1) ? and_ln890_1_fu_960_p2 : icmp_ln1019_3_fu_929_p2);

assign select_ln890_20_fu_5340_p3 = ((and_ln378_22_fu_5293_p2[0:0] == 1'b1) ? and_ln890_19_fu_5334_p2 : icmp_ln1019_41_fu_5303_p2);

assign select_ln890_21_fu_5583_p3 = ((and_ln378_23_fu_5536_p2[0:0] == 1'b1) ? and_ln890_20_fu_5577_p2 : icmp_ln1019_43_fu_5546_p2);

assign select_ln890_22_fu_5826_p3 = ((and_ln378_24_fu_5779_p2[0:0] == 1'b1) ? and_ln890_21_fu_5820_p2 : icmp_ln1019_45_fu_5789_p2);

assign select_ln890_23_fu_6056_p3 = ((and_ln378_25_fu_6009_p2[0:0] == 1'b1) ? and_ln890_22_fu_6050_p2 : icmp_ln1019_47_fu_6019_p2);

assign select_ln890_24_fu_6282_p3 = ((and_ln378_26_fu_6235_p2[0:0] == 1'b1) ? and_ln890_23_fu_6276_p2 : icmp_ln1019_49_fu_6245_p2);

assign select_ln890_3_fu_1209_p3 = ((and_ln378_3_fu_1162_p2[0:0] == 1'b1) ? and_ln890_2_fu_1203_p2 : icmp_ln1019_7_fu_1172_p2);

assign select_ln890_4_fu_1452_p3 = ((and_ln378_6_fu_1405_p2[0:0] == 1'b1) ? and_ln890_3_fu_1446_p2 : icmp_ln1019_9_fu_1415_p2);

assign select_ln890_5_fu_1695_p3 = ((and_ln378_7_fu_1648_p2[0:0] == 1'b1) ? and_ln890_4_fu_1689_p2 : icmp_ln1019_11_fu_1658_p2);

assign select_ln890_6_fu_1938_p3 = ((and_ln378_8_fu_1891_p2[0:0] == 1'b1) ? and_ln890_5_fu_1932_p2 : icmp_ln1019_13_fu_1901_p2);

assign select_ln890_7_fu_2181_p3 = ((and_ln378_9_fu_2134_p2[0:0] == 1'b1) ? and_ln890_6_fu_2175_p2 : icmp_ln1019_15_fu_2144_p2);

assign select_ln890_8_fu_2424_p3 = ((and_ln378_10_fu_2377_p2[0:0] == 1'b1) ? and_ln890_7_fu_2418_p2 : icmp_ln1019_17_fu_2387_p2);

assign select_ln890_9_fu_2667_p3 = ((and_ln378_11_fu_2620_p2[0:0] == 1'b1) ? and_ln890_8_fu_2661_p2 : icmp_ln1019_19_fu_2630_p2);

assign select_ln890_fu_723_p3 = ((and_ln378_fu_676_p2[0:0] == 1'b1) ? and_ln890_fu_717_p2 : icmp_ln1019_1_fu_686_p2);

assign sext_ln1273_10_cast_fu_442_p1 = $signed(sext_ln1273_10);

assign sext_ln1273_11_cast_fu_438_p1 = $signed(sext_ln1273_11);

assign sext_ln1273_12_cast_fu_434_p1 = $signed(sext_ln1273_12);

assign sext_ln1273_13_cast_fu_430_p1 = $signed(sext_ln1273_13);

assign sext_ln1273_14_cast_fu_426_p1 = $signed(sext_ln1273_14);

assign sext_ln1273_15_cast_fu_422_p1 = $signed(sext_ln1273_15);

assign sext_ln1273_16_cast_fu_418_p1 = $signed(sext_ln1273_16);

assign sext_ln1273_17_cast_fu_414_p1 = $signed(sext_ln1273_17);

assign sext_ln1273_18_cast_fu_410_p1 = $signed(sext_ln1273_18);

assign sext_ln1273_19_cast_fu_406_p1 = $signed(sext_ln1273_19);

assign sext_ln1273_1_cast_fu_478_p1 = $signed(sext_ln1273_1);

assign sext_ln1273_20_cast_fu_402_p1 = $signed(sext_ln1273_20);

assign sext_ln1273_21_cast_fu_398_p1 = $signed(sext_ln1273_21);

assign sext_ln1273_22_cast_fu_394_p1 = $signed(sext_ln1273_22);

assign sext_ln1273_23_cast_fu_390_p1 = $signed(sext_ln1273_23);

assign sext_ln1273_24_cast_fu_474_p1 = $signed(sext_ln1273_24);

assign sext_ln1273_3_cast_fu_470_p1 = $signed(sext_ln1273_3);

assign sext_ln1273_4_cast_fu_466_p1 = $signed(sext_ln1273_4);

assign sext_ln1273_5_cast_fu_462_p1 = $signed(sext_ln1273_5);

assign sext_ln1273_6_cast_fu_458_p1 = $signed(sext_ln1273_6);

assign sext_ln1273_7_cast_fu_454_p1 = $signed(sext_ln1273_7);

assign sext_ln1273_8_cast_fu_450_p1 = $signed(sext_ln1273_8);

assign sext_ln1273_9_cast_fu_446_p1 = $signed(sext_ln1273_9);

assign sext_ln1273_cast_fu_482_p1 = $signed(sext_ln1273);

assign sext_ln813_10_fu_2757_p1 = $signed(shl_ln838_5_fu_2749_p3);

assign sext_ln813_11_fu_3000_p1 = $signed(shl_ln838_7_fu_2992_p3);

assign sext_ln813_12_fu_3243_p1 = $signed(shl_ln838_8_fu_3235_p3);

assign sext_ln813_13_fu_3486_p1 = $signed(shl_ln838_10_fu_3478_p3);

assign sext_ln813_14_fu_3729_p1 = $signed(shl_ln838_11_fu_3721_p3);

assign sext_ln813_15_fu_3972_p1 = $signed(shl_ln838_12_fu_3964_p3);

assign sext_ln813_16_fu_4215_p1 = $signed(shl_ln838_13_fu_4207_p3);

assign sext_ln813_17_fu_4458_p1 = $signed(shl_ln838_14_fu_4450_p3);

assign sext_ln813_18_fu_4701_p1 = $signed(shl_ln838_15_fu_4693_p3);

assign sext_ln813_19_fu_4944_p1 = $signed(shl_ln838_16_fu_4936_p3);

assign sext_ln813_20_fu_5187_p1 = $signed(shl_ln838_17_fu_5179_p3);

assign sext_ln813_21_fu_5430_p1 = $signed(shl_ln838_18_fu_5422_p3);

assign sext_ln813_22_fu_5673_p1 = $signed(shl_ln838_19_fu_5665_p3);

assign sext_ln813_23_fu_5916_p1 = $signed(shl_ln838_20_fu_5908_p3);

assign sext_ln813_24_fu_6146_p1 = $signed(shl_ln838_21_fu_6138_p3);

assign sext_ln813_3_fu_813_p1 = $signed(shl_ln_fu_805_p3);

assign sext_ln813_4_fu_1056_p1 = $signed(shl_ln838_1_fu_1048_p3);

assign sext_ln813_5_fu_1299_p1 = $signed(shl_ln838_3_fu_1291_p3);

assign sext_ln813_6_fu_1542_p1 = $signed(shl_ln838_6_fu_1534_p3);

assign sext_ln813_7_fu_1785_p1 = $signed(shl_ln838_9_fu_1777_p3);

assign sext_ln813_8_fu_2028_p1 = $signed(shl_ln838_s_fu_2020_p3);

assign sext_ln813_9_fu_2514_p1 = $signed(shl_ln838_4_fu_2506_p3);

assign sext_ln813_fu_2271_p1 = $signed(shl_ln838_2_fu_2263_p3);

assign shl_ln838_10_fu_3478_p3 = {{select_ln346_24_fu_3470_p3}, {16'd0}};

assign shl_ln838_11_fu_3721_p3 = {{select_ln346_26_fu_3713_p3}, {16'd0}};

assign shl_ln838_12_fu_3964_p3 = {{select_ln346_28_fu_3956_p3}, {16'd0}};

assign shl_ln838_13_fu_4207_p3 = {{select_ln346_30_fu_4199_p3}, {16'd0}};

assign shl_ln838_14_fu_4450_p3 = {{select_ln346_32_fu_4442_p3}, {16'd0}};

assign shl_ln838_15_fu_4693_p3 = {{select_ln346_34_fu_4685_p3}, {16'd0}};

assign shl_ln838_16_fu_4936_p3 = {{select_ln346_36_fu_4928_p3}, {16'd0}};

assign shl_ln838_17_fu_5179_p3 = {{select_ln346_38_fu_5171_p3}, {16'd0}};

assign shl_ln838_18_fu_5422_p3 = {{select_ln346_40_fu_5414_p3}, {16'd0}};

assign shl_ln838_19_fu_5665_p3 = {{select_ln346_42_fu_5657_p3}, {16'd0}};

assign shl_ln838_1_fu_1048_p3 = {{select_ln346_5_fu_1040_p3}, {16'd0}};

assign shl_ln838_20_fu_5908_p3 = {{select_ln346_44_fu_5900_p3}, {16'd0}};

assign shl_ln838_21_fu_6138_p3 = {{select_ln346_46_fu_6130_p3}, {16'd0}};

assign shl_ln838_2_fu_2263_p3 = {{select_ln346_fu_2255_p3}, {16'd0}};

assign shl_ln838_3_fu_1291_p3 = {{select_ln346_7_fu_1283_p3}, {16'd0}};

assign shl_ln838_4_fu_2506_p3 = {{select_ln346_16_fu_2498_p3}, {16'd0}};

assign shl_ln838_5_fu_2749_p3 = {{select_ln346_18_fu_2741_p3}, {16'd0}};

assign shl_ln838_6_fu_1534_p3 = {{select_ln346_9_fu_1526_p3}, {16'd0}};

assign shl_ln838_7_fu_2992_p3 = {{select_ln346_20_fu_2984_p3}, {16'd0}};

assign shl_ln838_8_fu_3235_p3 = {{select_ln346_22_fu_3227_p3}, {16'd0}};

assign shl_ln838_9_fu_1777_p3 = {{select_ln346_11_fu_1769_p3}, {16'd0}};

assign shl_ln838_s_fu_2020_p3 = {{select_ln346_13_fu_2012_p3}, {16'd0}};

assign shl_ln_fu_805_p3 = {{select_ln346_3_fu_797_p3}, {16'd0}};

assign temp1_V_0_1_out = temp1_V_3_2_fu_178;

assign temp1_V_1_1_out = temp1_V_3_3_fu_182;

assign temp1_V_2_1_out = temp1_V_3_4_fu_186;

assign temp1_V_3_1_out = temp1_V_3_1_fu_190;

assign temp1_V_3_6_fu_6399_p3 = ((icmp_ln1420_2_fu_6374_p2[0:0] == 1'b1) ? temp1_V_3_9_fu_6356_p3 : temp1_V_3_4_fu_186);

assign temp1_V_3_7_fu_6407_p3 = ((icmp_ln1420_1_fu_6369_p2[0:0] == 1'b1) ? temp1_V_3_9_fu_6356_p3 : temp1_V_3_3_fu_182);

assign temp1_V_3_8_fu_6415_p3 = ((icmp_ln1420_fu_6364_p2[0:0] == 1'b1) ? temp1_V_3_9_fu_6356_p3 : temp1_V_3_2_fu_178);

assign temp1_V_3_9_fu_6356_p3 = ((or_ln346_26_fu_6350_p2[0:0] == 1'b1) ? select_ln346_47_fu_6342_p3 : add_ln377_26_fu_6216_p2);

assign temp1_V_3_fu_6391_p3 = ((or_ln1420_1_fu_6385_p2[0:0] == 1'b1) ? temp1_V_3_1_fu_190 : temp1_V_3_9_fu_6356_p3);

assign tmp_101_fu_1877_p3 = add_ln377_8_fu_1872_p2[32'd31];

assign tmp_102_fu_1919_p3 = add_ln1347_5_reg_6901[32'd48];

assign tmp_106_fu_2120_p3 = add_ln377_9_fu_2115_p2[32'd31];

assign tmp_107_fu_2162_p3 = add_ln1347_6_reg_6948[32'd48];

assign tmp_111_fu_2363_p3 = add_ln377_10_fu_2358_p2[32'd31];

assign tmp_112_fu_2405_p3 = add_ln1347_7_reg_6995[32'd48];

assign tmp_116_fu_2606_p3 = add_ln377_11_fu_2601_p2[32'd31];

assign tmp_117_fu_2648_p3 = add_ln1347_8_reg_7042[32'd48];

assign tmp_121_fu_2849_p3 = add_ln377_12_fu_2844_p2[32'd31];

assign tmp_122_fu_2891_p3 = add_ln1347_9_reg_7089[32'd48];

assign tmp_126_fu_3092_p3 = add_ln377_13_fu_3087_p2[32'd31];

assign tmp_127_fu_3134_p3 = add_ln1347_10_reg_7136[32'd48];

assign tmp_131_fu_3335_p3 = add_ln377_14_fu_3330_p2[32'd31];

assign tmp_132_fu_3377_p3 = add_ln1347_11_reg_7183[32'd48];

assign tmp_136_fu_3578_p3 = add_ln377_15_fu_3573_p2[32'd31];

assign tmp_137_fu_3620_p3 = add_ln1347_12_reg_7230[32'd48];

assign tmp_141_fu_3821_p3 = add_ln377_16_fu_3816_p2[32'd31];

assign tmp_142_fu_3863_p3 = add_ln1347_13_reg_7277[32'd48];

assign tmp_146_fu_4064_p3 = add_ln377_17_fu_4059_p2[32'd31];

assign tmp_147_fu_4106_p3 = add_ln1347_14_reg_7324[32'd48];

assign tmp_151_fu_4307_p3 = add_ln377_18_fu_4302_p2[32'd31];

assign tmp_152_fu_4349_p3 = add_ln1347_15_reg_7371[32'd48];

assign tmp_156_fu_4550_p3 = add_ln377_19_fu_4545_p2[32'd31];

assign tmp_157_fu_4592_p3 = add_ln1347_16_reg_7418[32'd48];

assign tmp_161_fu_4793_p3 = add_ln377_20_fu_4788_p2[32'd31];

assign tmp_162_fu_4835_p3 = add_ln1347_17_reg_7465[32'd48];

assign tmp_166_fu_5036_p3 = add_ln377_21_fu_5031_p2[32'd31];

assign tmp_167_fu_5078_p3 = add_ln1347_18_reg_7512[32'd48];

assign tmp_171_fu_5279_p3 = add_ln377_22_fu_5274_p2[32'd31];

assign tmp_172_fu_5321_p3 = add_ln1347_19_reg_7559[32'd48];

assign tmp_176_fu_5522_p3 = add_ln377_23_fu_5517_p2[32'd31];

assign tmp_177_fu_5564_p3 = add_ln1347_20_reg_7606[32'd48];

assign tmp_181_fu_5765_p3 = add_ln377_24_fu_5760_p2[32'd31];

assign tmp_182_fu_5807_p3 = add_ln1347_21_reg_7653[32'd48];

assign tmp_186_fu_5995_p3 = add_ln377_25_fu_5990_p2[32'd31];

assign tmp_187_fu_6037_p3 = add_ln1347_22_reg_7700[32'd48];

assign tmp_191_fu_6221_p3 = add_ln377_26_fu_6216_p2[32'd31];

assign tmp_192_fu_6263_p3 = add_ln1347_23_reg_7742[32'd48];

assign tmp_76_fu_662_p3 = add_ln377_fu_657_p2[32'd31];

assign tmp_77_fu_704_p3 = mul_ln1273_reg_6661[32'd48];

assign tmp_81_fu_905_p3 = add_ln377_1_fu_900_p2[32'd31];

assign tmp_82_fu_947_p3 = add_ln1347_reg_6713[32'd48];

assign tmp_86_fu_1148_p3 = add_ln377_3_fu_1143_p2[32'd31];

assign tmp_87_fu_1190_p3 = add_ln1347_1_reg_6760[32'd48];

assign tmp_91_fu_1391_p3 = add_ln377_6_fu_1386_p2[32'd31];

assign tmp_92_fu_1433_p3 = add_ln1347_3_reg_6807[32'd48];

assign tmp_96_fu_1634_p3 = add_ln377_7_fu_1629_p2[32'd31];

assign tmp_97_fu_1676_p3 = add_ln1347_4_reg_6854[32'd48];

assign trunc_ln25_fu_526_p1 = ap_sig_allocacmp_i[1:0];

assign xor_ln890_10_fu_1683_p2 = (tmp_97_fu_1676_p3 ^ 1'd1);

assign xor_ln890_11_fu_1926_p2 = (tmp_102_fu_1919_p3 ^ 1'd1);

assign xor_ln890_12_fu_2169_p2 = (tmp_107_fu_2162_p3 ^ 1'd1);

assign xor_ln890_13_fu_2412_p2 = (tmp_112_fu_2405_p3 ^ 1'd1);

assign xor_ln890_14_fu_2655_p2 = (tmp_117_fu_2648_p3 ^ 1'd1);

assign xor_ln890_15_fu_2898_p2 = (tmp_122_fu_2891_p3 ^ 1'd1);

assign xor_ln890_16_fu_3141_p2 = (tmp_127_fu_3134_p3 ^ 1'd1);

assign xor_ln890_17_fu_3384_p2 = (tmp_132_fu_3377_p3 ^ 1'd1);

assign xor_ln890_18_fu_3627_p2 = (tmp_137_fu_3620_p3 ^ 1'd1);

assign xor_ln890_19_fu_3870_p2 = (tmp_142_fu_3863_p3 ^ 1'd1);

assign xor_ln890_20_fu_4113_p2 = (tmp_147_fu_4106_p3 ^ 1'd1);

assign xor_ln890_21_fu_4356_p2 = (tmp_152_fu_4349_p3 ^ 1'd1);

assign xor_ln890_22_fu_4599_p2 = (tmp_157_fu_4592_p3 ^ 1'd1);

assign xor_ln890_23_fu_4842_p2 = (tmp_162_fu_4835_p3 ^ 1'd1);

assign xor_ln890_24_fu_5085_p2 = (tmp_167_fu_5078_p3 ^ 1'd1);

assign xor_ln890_25_fu_5328_p2 = (tmp_172_fu_5321_p3 ^ 1'd1);

assign xor_ln890_26_fu_5571_p2 = (tmp_177_fu_5564_p3 ^ 1'd1);

assign xor_ln890_27_fu_5814_p2 = (tmp_182_fu_5807_p3 ^ 1'd1);

assign xor_ln890_28_fu_6044_p2 = (tmp_187_fu_6037_p3 ^ 1'd1);

assign xor_ln890_29_fu_6270_p2 = (tmp_192_fu_6263_p3 ^ 1'd1);

assign xor_ln890_7_fu_954_p2 = (tmp_82_fu_947_p3 ^ 1'd1);

assign xor_ln890_8_fu_1197_p2 = (tmp_87_fu_1190_p3 ^ 1'd1);

assign xor_ln890_9_fu_1440_p2 = (tmp_92_fu_1433_p3 ^ 1'd1);

assign xor_ln890_fu_711_p2 = (tmp_77_fu_704_p3 ^ 1'd1);

assign xor_ln895_10_fu_1223_p2 = (select_ln888_3_fu_1182_p3 ^ 1'd1);

assign xor_ln895_11_fu_1235_p2 = (tmp_83_reg_6765 ^ 1'd1);

assign xor_ln895_14_fu_1478_p2 = (tmp_88_reg_6812 ^ 1'd1);

assign xor_ln895_15_fu_1709_p2 = (select_ln888_5_fu_1668_p3 ^ 1'd1);

assign xor_ln895_16_fu_1721_p2 = (tmp_93_reg_6859 ^ 1'd1);

assign xor_ln895_17_fu_1952_p2 = (select_ln888_6_fu_1911_p3 ^ 1'd1);

assign xor_ln895_18_fu_1964_p2 = (tmp_98_reg_6906 ^ 1'd1);

assign xor_ln895_19_fu_2195_p2 = (select_ln888_7_fu_2154_p3 ^ 1'd1);

assign xor_ln895_20_fu_2207_p2 = (tmp_103_reg_6953 ^ 1'd1);

assign xor_ln895_21_fu_2438_p2 = (select_ln888_8_fu_2397_p3 ^ 1'd1);

assign xor_ln895_22_fu_2450_p2 = (tmp_108_reg_7000 ^ 1'd1);

assign xor_ln895_23_fu_2681_p2 = (select_ln888_9_fu_2640_p3 ^ 1'd1);

assign xor_ln895_24_fu_2693_p2 = (tmp_113_reg_7047 ^ 1'd1);

assign xor_ln895_25_fu_2924_p2 = (select_ln888_10_fu_2883_p3 ^ 1'd1);

assign xor_ln895_26_fu_2936_p2 = (tmp_118_reg_7094 ^ 1'd1);

assign xor_ln895_27_fu_3167_p2 = (select_ln888_11_fu_3126_p3 ^ 1'd1);

assign xor_ln895_28_fu_3179_p2 = (tmp_123_reg_7141 ^ 1'd1);

assign xor_ln895_29_fu_3410_p2 = (select_ln888_12_fu_3369_p3 ^ 1'd1);

assign xor_ln895_2_fu_737_p2 = (select_ln888_fu_696_p3 ^ 1'd1);

assign xor_ln895_30_fu_3422_p2 = (tmp_128_reg_7188 ^ 1'd1);

assign xor_ln895_31_fu_3653_p2 = (select_ln888_13_fu_3612_p3 ^ 1'd1);

assign xor_ln895_32_fu_3665_p2 = (tmp_133_reg_7235 ^ 1'd1);

assign xor_ln895_33_fu_3896_p2 = (select_ln888_14_fu_3855_p3 ^ 1'd1);

assign xor_ln895_34_fu_3908_p2 = (tmp_138_reg_7282 ^ 1'd1);

assign xor_ln895_35_fu_4139_p2 = (select_ln888_15_fu_4098_p3 ^ 1'd1);

assign xor_ln895_36_fu_4151_p2 = (tmp_143_reg_7329 ^ 1'd1);

assign xor_ln895_37_fu_4382_p2 = (select_ln888_16_fu_4341_p3 ^ 1'd1);

assign xor_ln895_38_fu_4394_p2 = (tmp_148_reg_7376 ^ 1'd1);

assign xor_ln895_39_fu_4625_p2 = (select_ln888_17_fu_4584_p3 ^ 1'd1);

assign xor_ln895_3_fu_749_p2 = (tmp_73_reg_6666 ^ 1'd1);

assign xor_ln895_40_fu_4637_p2 = (tmp_153_reg_7423 ^ 1'd1);

assign xor_ln895_41_fu_4868_p2 = (select_ln888_18_fu_4827_p3 ^ 1'd1);

assign xor_ln895_42_fu_4880_p2 = (tmp_158_reg_7470 ^ 1'd1);

assign xor_ln895_43_fu_5111_p2 = (select_ln888_19_fu_5070_p3 ^ 1'd1);

assign xor_ln895_44_fu_5123_p2 = (tmp_163_reg_7517 ^ 1'd1);

assign xor_ln895_45_fu_5354_p2 = (select_ln888_20_fu_5313_p3 ^ 1'd1);

assign xor_ln895_46_fu_5366_p2 = (tmp_168_reg_7564 ^ 1'd1);

assign xor_ln895_47_fu_5597_p2 = (select_ln888_21_fu_5556_p3 ^ 1'd1);

assign xor_ln895_48_fu_5609_p2 = (tmp_173_reg_7611 ^ 1'd1);

assign xor_ln895_49_fu_5840_p2 = (select_ln888_22_fu_5799_p3 ^ 1'd1);

assign xor_ln895_4_fu_980_p2 = (select_ln888_1_fu_939_p3 ^ 1'd1);

assign xor_ln895_50_fu_5852_p2 = (tmp_178_reg_7658 ^ 1'd1);

assign xor_ln895_51_fu_6070_p2 = (select_ln888_23_fu_6029_p3 ^ 1'd1);

assign xor_ln895_52_fu_6082_p2 = (tmp_183_reg_7705 ^ 1'd1);

assign xor_ln895_53_fu_6296_p2 = (select_ln888_24_fu_6255_p3 ^ 1'd1);

assign xor_ln895_54_fu_6308_p2 = (tmp_188_reg_7747 ^ 1'd1);

assign xor_ln895_5_fu_992_p2 = (tmp_78_reg_6718 ^ 1'd1);

assign xor_ln895_fu_1466_p2 = (select_ln888_4_fu_1425_p3 ^ 1'd1);

assign xor_ln896_10_fu_1399_p2 = (tmp_91_fu_1391_p3 ^ 1'd1);

assign xor_ln896_15_fu_1489_p2 = (select_ln890_4_fu_1452_p3 ^ 1'd1);

assign xor_ln896_16_fu_1642_p2 = (tmp_96_fu_1634_p3 ^ 1'd1);

assign xor_ln896_1_fu_760_p2 = (select_ln890_fu_723_p3 ^ 1'd1);

assign xor_ln896_20_fu_772_p2 = (or_ln896_fu_766_p2 ^ and_ln891_fu_731_p2);

assign xor_ln896_21_fu_1732_p2 = (select_ln890_5_fu_1695_p3 ^ 1'd1);

assign xor_ln896_22_fu_1885_p2 = (tmp_101_fu_1877_p3 ^ 1'd1);

assign xor_ln896_23_fu_1015_p2 = (or_ln896_1_fu_1009_p2 ^ and_ln891_1_fu_974_p2);

assign xor_ln896_24_fu_1258_p2 = (or_ln896_18_fu_1252_p2 ^ and_ln891_24_fu_1217_p2);

assign xor_ln896_25_fu_1501_p2 = (or_ln896_3_fu_1495_p2 ^ and_ln891_3_fu_1460_p2);

assign xor_ln896_26_fu_1975_p2 = (select_ln890_6_fu_1938_p3 ^ 1'd1);

assign xor_ln896_27_fu_2128_p2 = (tmp_106_fu_2120_p3 ^ 1'd1);

assign xor_ln896_28_fu_1744_p2 = (or_ln896_4_fu_1738_p2 ^ and_ln891_4_fu_1703_p2);

assign xor_ln896_29_fu_2218_p2 = (select_ln890_7_fu_2181_p3 ^ 1'd1);

assign xor_ln896_2_fu_913_p2 = (tmp_81_fu_905_p3 ^ 1'd1);

assign xor_ln896_30_fu_2371_p2 = (tmp_111_fu_2363_p3 ^ 1'd1);

assign xor_ln896_31_fu_2461_p2 = (select_ln890_8_fu_2424_p3 ^ 1'd1);

assign xor_ln896_32_fu_2614_p2 = (tmp_116_fu_2606_p3 ^ 1'd1);

assign xor_ln896_33_fu_2704_p2 = (select_ln890_9_fu_2667_p3 ^ 1'd1);

assign xor_ln896_34_fu_2857_p2 = (tmp_121_fu_2849_p3 ^ 1'd1);

assign xor_ln896_35_fu_2947_p2 = (select_ln890_10_fu_2910_p3 ^ 1'd1);

assign xor_ln896_36_fu_3100_p2 = (tmp_126_fu_3092_p3 ^ 1'd1);

assign xor_ln896_37_fu_3190_p2 = (select_ln890_11_fu_3153_p3 ^ 1'd1);

assign xor_ln896_38_fu_3343_p2 = (tmp_131_fu_3335_p3 ^ 1'd1);

assign xor_ln896_39_fu_3433_p2 = (select_ln890_12_fu_3396_p3 ^ 1'd1);

assign xor_ln896_40_fu_3586_p2 = (tmp_136_fu_3578_p3 ^ 1'd1);

assign xor_ln896_41_fu_3676_p2 = (select_ln890_13_fu_3639_p3 ^ 1'd1);

assign xor_ln896_42_fu_3829_p2 = (tmp_141_fu_3821_p3 ^ 1'd1);

assign xor_ln896_43_fu_3919_p2 = (select_ln890_14_fu_3882_p3 ^ 1'd1);

assign xor_ln896_44_fu_4072_p2 = (tmp_146_fu_4064_p3 ^ 1'd1);

assign xor_ln896_45_fu_4162_p2 = (select_ln890_15_fu_4125_p3 ^ 1'd1);

assign xor_ln896_46_fu_4315_p2 = (tmp_151_fu_4307_p3 ^ 1'd1);

assign xor_ln896_47_fu_4405_p2 = (select_ln890_16_fu_4368_p3 ^ 1'd1);

assign xor_ln896_48_fu_4558_p2 = (tmp_156_fu_4550_p3 ^ 1'd1);

assign xor_ln896_49_fu_4648_p2 = (select_ln890_17_fu_4611_p3 ^ 1'd1);

assign xor_ln896_4_fu_1003_p2 = (select_ln890_1_fu_966_p3 ^ 1'd1);

assign xor_ln896_50_fu_4801_p2 = (tmp_161_fu_4793_p3 ^ 1'd1);

assign xor_ln896_51_fu_4891_p2 = (select_ln890_18_fu_4854_p3 ^ 1'd1);

assign xor_ln896_52_fu_5044_p2 = (tmp_166_fu_5036_p3 ^ 1'd1);

assign xor_ln896_53_fu_5134_p2 = (select_ln890_19_fu_5097_p3 ^ 1'd1);

assign xor_ln896_54_fu_5287_p2 = (tmp_171_fu_5279_p3 ^ 1'd1);

assign xor_ln896_55_fu_5377_p2 = (select_ln890_20_fu_5340_p3 ^ 1'd1);

assign xor_ln896_56_fu_5530_p2 = (tmp_176_fu_5522_p3 ^ 1'd1);

assign xor_ln896_57_fu_5620_p2 = (select_ln890_21_fu_5583_p3 ^ 1'd1);

assign xor_ln896_58_fu_5773_p2 = (tmp_181_fu_5765_p3 ^ 1'd1);

assign xor_ln896_59_fu_5863_p2 = (select_ln890_22_fu_5826_p3 ^ 1'd1);

assign xor_ln896_5_fu_1156_p2 = (tmp_86_fu_1148_p3 ^ 1'd1);

assign xor_ln896_60_fu_6003_p2 = (tmp_186_fu_5995_p3 ^ 1'd1);

assign xor_ln896_61_fu_6093_p2 = (select_ln890_23_fu_6056_p3 ^ 1'd1);

assign xor_ln896_62_fu_6229_p2 = (tmp_191_fu_6221_p3 ^ 1'd1);

assign xor_ln896_63_fu_6319_p2 = (select_ln890_24_fu_6282_p3 ^ 1'd1);

assign xor_ln896_64_fu_1987_p2 = (or_ln896_5_fu_1981_p2 ^ and_ln891_5_fu_1946_p2);

assign xor_ln896_65_fu_2230_p2 = (or_ln896_6_fu_2224_p2 ^ and_ln891_6_fu_2189_p2);

assign xor_ln896_66_fu_2473_p2 = (or_ln896_7_fu_2467_p2 ^ and_ln891_7_fu_2432_p2);

assign xor_ln896_67_fu_2716_p2 = (or_ln896_8_fu_2710_p2 ^ and_ln891_8_fu_2675_p2);

assign xor_ln896_68_fu_2959_p2 = (or_ln896_9_fu_2953_p2 ^ and_ln891_9_fu_2918_p2);

assign xor_ln896_69_fu_3202_p2 = (or_ln896_10_fu_3196_p2 ^ and_ln891_10_fu_3161_p2);

assign xor_ln896_70_fu_3445_p2 = (or_ln896_11_fu_3439_p2 ^ and_ln891_11_fu_3404_p2);

assign xor_ln896_71_fu_3688_p2 = (or_ln896_12_fu_3682_p2 ^ and_ln891_12_fu_3647_p2);

assign xor_ln896_72_fu_3931_p2 = (or_ln896_13_fu_3925_p2 ^ and_ln891_13_fu_3890_p2);

assign xor_ln896_73_fu_4174_p2 = (or_ln896_14_fu_4168_p2 ^ and_ln891_14_fu_4133_p2);

assign xor_ln896_74_fu_4417_p2 = (or_ln896_15_fu_4411_p2 ^ and_ln891_15_fu_4376_p2);

assign xor_ln896_75_fu_4660_p2 = (or_ln896_16_fu_4654_p2 ^ and_ln891_16_fu_4619_p2);

assign xor_ln896_76_fu_4903_p2 = (or_ln896_17_fu_4897_p2 ^ and_ln891_17_fu_4862_p2);

assign xor_ln896_77_fu_5146_p2 = (or_ln896_24_fu_5140_p2 ^ and_ln891_18_fu_5105_p2);

assign xor_ln896_78_fu_5389_p2 = (or_ln896_19_fu_5383_p2 ^ and_ln891_19_fu_5348_p2);

assign xor_ln896_79_fu_5632_p2 = (or_ln896_20_fu_5626_p2 ^ and_ln891_20_fu_5591_p2);

assign xor_ln896_80_fu_5875_p2 = (or_ln896_21_fu_5869_p2 ^ and_ln891_21_fu_5834_p2);

assign xor_ln896_81_fu_6105_p2 = (or_ln896_22_fu_6099_p2 ^ and_ln891_22_fu_6064_p2);

assign xor_ln896_82_fu_6331_p2 = (or_ln896_23_fu_6325_p2 ^ and_ln891_23_fu_6290_p2);

assign xor_ln896_9_fu_1246_p2 = (select_ln890_3_fu_1209_p3 ^ 1'd1);

assign xor_ln896_fu_670_p2 = (tmp_76_fu_662_p3 ^ 1'd1);

assign zext_ln377_10_fu_3084_p1 = tmp_125_reg_7126_pp0_iter11_reg;

assign zext_ln377_11_fu_3327_p1 = tmp_130_reg_7173_pp0_iter12_reg;

assign zext_ln377_12_fu_3570_p1 = tmp_135_reg_7220_pp0_iter13_reg;

assign zext_ln377_13_fu_3813_p1 = tmp_140_reg_7267_pp0_iter14_reg;

assign zext_ln377_14_fu_4056_p1 = tmp_145_reg_7314_pp0_iter15_reg;

assign zext_ln377_15_fu_4299_p1 = tmp_150_reg_7361_pp0_iter16_reg;

assign zext_ln377_16_fu_4542_p1 = tmp_155_reg_7408_pp0_iter17_reg;

assign zext_ln377_17_fu_4785_p1 = tmp_160_reg_7455_pp0_iter18_reg;

assign zext_ln377_18_fu_5028_p1 = tmp_165_reg_7502_pp0_iter19_reg;

assign zext_ln377_19_fu_5271_p1 = tmp_170_reg_7549_pp0_iter20_reg;

assign zext_ln377_1_fu_897_p1 = tmp_80_reg_6703_pp0_iter2_reg;

assign zext_ln377_20_fu_5514_p1 = tmp_175_reg_7596_pp0_iter21_reg;

assign zext_ln377_21_fu_5757_p1 = tmp_180_reg_7643_pp0_iter22_reg;

assign zext_ln377_22_fu_5987_p1 = tmp_185_reg_7690_pp0_iter23_reg;

assign zext_ln377_23_fu_6213_p1 = tmp_190_reg_7737_pp0_iter24_reg;

assign zext_ln377_2_fu_1140_p1 = tmp_85_reg_6750_pp0_iter3_reg;

assign zext_ln377_3_fu_1383_p1 = tmp_90_reg_6797_pp0_iter4_reg;

assign zext_ln377_4_fu_1626_p1 = tmp_95_reg_6844_pp0_iter5_reg;

assign zext_ln377_5_fu_1869_p1 = tmp_100_reg_6891_pp0_iter6_reg;

assign zext_ln377_6_fu_2112_p1 = tmp_105_reg_6938_pp0_iter7_reg;

assign zext_ln377_7_fu_2355_p1 = tmp_110_reg_6985_pp0_iter8_reg;

assign zext_ln377_8_fu_2598_p1 = tmp_115_reg_7032_pp0_iter9_reg;

assign zext_ln377_9_fu_2841_p1 = tmp_120_reg_7079_pp0_iter10_reg;

assign zext_ln377_fu_654_p1 = tmp_75_reg_6682;

endmodule //mpc_qp_admm_Pipeline_mvmult_row
