module motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config5_s (
        ap_clk,
        ap_rst,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [31:0] p_read;
input  [31:0] p_read1;
input  [31:0] p_read2;
input  [31:0] p_read3;
input  [31:0] p_read4;
input  [31:0] p_read5;
input  [31:0] p_read6;
input  [31:0] p_read7;
input  [31:0] p_read8;
output  [31:0] ap_return_0;
output  [31:0] ap_return_1;
output  [31:0] ap_return_2;
output  [31:0] ap_return_3;
output  [31:0] ap_return_4;
output  [31:0] ap_return_5;
output  [31:0] ap_return_6;
output  [31:0] ap_return_7;
output  [31:0] ap_return_8;
input   ap_ce;

reg[31:0] ap_return_0;
reg[31:0] ap_return_1;
reg[31:0] ap_return_2;
reg[31:0] ap_return_3;
reg[31:0] ap_return_4;
reg[31:0] ap_return_5;
reg[31:0] ap_return_6;
reg[31:0] ap_return_7;
reg[31:0] ap_return_8;

wire   [41:0] r_V_fu_536_p2;
reg   [41:0] r_V_reg_9071;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [42:0] r_V_78_fu_527_p2;
reg   [42:0] r_V_78_reg_9075;
wire   [43:0] r_V_79_fu_484_p2;
reg   [43:0] r_V_79_reg_9079;
wire   [41:0] r_V_80_fu_509_p2;
reg   [41:0] r_V_80_reg_9083;
wire   [41:0] r_V_81_fu_489_p2;
reg   [41:0] r_V_81_reg_9087;
wire   [43:0] r_V_82_fu_497_p2;
reg   [43:0] r_V_82_reg_9091;
wire   [44:0] r_V_83_fu_507_p2;
reg   [44:0] r_V_83_reg_9095;
wire   [39:0] r_V_84_fu_494_p2;
reg   [39:0] r_V_84_reg_9099;
wire   [42:0] r_V_85_fu_495_p2;
reg   [42:0] r_V_85_reg_9103;
wire   [44:0] r_V_86_fu_505_p2;
reg   [44:0] r_V_86_reg_9107;
wire   [41:0] r_V_87_fu_538_p2;
reg   [41:0] r_V_87_reg_9111;
wire   [39:0] r_V_88_fu_498_p2;
reg   [39:0] r_V_88_reg_9115;
wire   [43:0] r_V_89_fu_482_p2;
reg   [43:0] r_V_89_reg_9119;
wire   [41:0] r_V_90_fu_480_p2;
reg   [41:0] r_V_90_reg_9123;
wire   [41:0] r_V_92_fu_522_p2;
reg   [41:0] r_V_92_reg_9127;
wire   [42:0] r_V_93_fu_532_p2;
reg   [42:0] r_V_93_reg_9131;
wire   [38:0] r_V_94_fu_499_p2;
reg   [38:0] r_V_94_reg_9135;
wire   [54:0] r_V_95_fu_503_p2;
reg   [54:0] r_V_95_reg_9139;
wire   [43:0] r_V_96_fu_530_p2;
reg   [43:0] r_V_96_reg_9143;
wire   [40:0] r_V_97_fu_504_p2;
reg   [40:0] r_V_97_reg_9147;
wire   [55:0] r_V_98_fu_501_p2;
reg   [55:0] r_V_98_reg_9151;
wire   [51:0] r_V_99_fu_465_p2;
reg   [51:0] r_V_99_reg_9155;
wire   [44:0] r_V_100_fu_534_p2;
reg   [44:0] r_V_100_reg_9159;
wire   [42:0] r_V_101_fu_478_p2;
reg   [42:0] r_V_101_reg_9163;
wire   [40:0] r_V_102_fu_474_p2;
reg   [40:0] r_V_102_reg_9167;
wire   [46:0] r_V_103_fu_469_p2;
reg   [46:0] r_V_103_reg_9171;
wire   [41:0] r_V_104_fu_466_p2;
reg   [41:0] r_V_104_reg_12983;
wire   [42:0] r_V_105_fu_539_p2;
reg   [42:0] r_V_105_reg_12987;
wire   [41:0] r_V_106_fu_512_p2;
reg   [41:0] r_V_106_reg_12991;
wire   [42:0] r_V_107_fu_463_p2;
reg   [42:0] r_V_107_reg_12995;
wire   [43:0] r_V_108_fu_529_p2;
reg   [43:0] r_V_108_reg_12999;
wire   [41:0] r_V_109_fu_485_p2;
reg   [41:0] r_V_109_reg_13003;
wire   [43:0] r_V_111_fu_526_p2;
reg   [43:0] r_V_111_reg_13007;
wire   [42:0] r_V_112_fu_471_p2;
reg   [42:0] r_V_112_reg_13011;
wire   [54:0] r_V_113_fu_535_p2;
reg   [54:0] r_V_113_reg_13015;
wire   [41:0] r_V_114_fu_475_p2;
reg   [41:0] r_V_114_reg_13019;
wire   [44:0] r_V_115_fu_468_p2;
reg   [44:0] r_V_115_reg_13023;
wire   [44:0] r_V_116_fu_537_p2;
reg   [44:0] r_V_116_reg_13027;
wire   [46:0] r_V_117_fu_519_p2;
reg   [46:0] r_V_117_reg_13031;
wire   [42:0] r_V_118_fu_470_p2;
reg   [42:0] r_V_118_reg_13035;
wire   [44:0] r_V_119_fu_542_p2;
reg   [44:0] r_V_119_reg_13039;
wire   [43:0] r_V_120_fu_520_p2;
reg   [43:0] r_V_120_reg_13043;
wire   [43:0] r_V_121_fu_477_p2;
reg   [43:0] r_V_121_reg_13047;
wire   [42:0] r_V_123_fu_472_p2;
reg   [42:0] r_V_123_reg_15547;
wire   [43:0] r_V_124_fu_462_p2;
reg   [43:0] r_V_124_reg_15551;
wire   [42:0] r_V_125_fu_510_p2;
reg   [42:0] r_V_125_reg_15555;
wire   [43:0] r_V_126_fu_515_p2;
reg   [43:0] r_V_126_reg_15559;
wire   [42:0] r_V_127_fu_479_p2;
reg   [42:0] r_V_127_reg_15563;
wire   [44:0] r_V_128_fu_513_p2;
reg   [44:0] r_V_128_reg_15567;
wire   [39:0] r_V_129_fu_521_p2;
reg   [39:0] r_V_129_reg_15571;
wire   [41:0] r_V_130_fu_491_p2;
reg   [41:0] r_V_130_reg_15575;
wire   [43:0] r_V_131_fu_506_p2;
reg   [43:0] r_V_131_reg_15579;
wire   [42:0] r_V_132_fu_533_p2;
reg   [42:0] r_V_132_reg_15583;
wire   [42:0] r_V_133_fu_486_p2;
reg   [42:0] r_V_133_reg_15587;
wire   [43:0] r_V_134_fu_525_p2;
reg   [43:0] r_V_134_reg_15591;
wire   [42:0] r_V_135_fu_496_p2;
reg   [42:0] r_V_135_reg_15595;
wire   [42:0] r_V_136_fu_500_p2;
reg   [42:0] r_V_136_reg_15599;
wire   [40:0] r_V_137_fu_464_p2;
reg   [40:0] r_V_137_reg_15603;
wire   [41:0] r_V_138_fu_528_p2;
reg   [41:0] r_V_138_reg_15607;
wire   [54:0] r_V_140_fu_481_p2;
reg   [54:0] r_V_140_reg_17175;
wire   [43:0] r_V_141_fu_541_p2;
reg   [43:0] r_V_141_reg_17179;
wire   [42:0] r_V_142_fu_492_p2;
reg   [42:0] r_V_142_reg_17183;
wire   [49:0] r_V_143_fu_540_p2;
reg   [49:0] r_V_143_reg_17187;
wire   [48:0] r_V_144_fu_490_p2;
reg   [48:0] r_V_144_reg_17191;
wire   [43:0] r_V_145_fu_476_p2;
reg   [43:0] r_V_145_reg_17195;
wire   [43:0] r_V_146_fu_514_p2;
reg   [43:0] r_V_146_reg_17199;
wire   [43:0] r_V_147_fu_508_p2;
reg   [43:0] r_V_147_reg_17203;
wire   [48:0] r_V_148_fu_518_p2;
reg   [48:0] r_V_148_reg_17207;
wire   [54:0] r_V_149_fu_493_p2;
reg   [54:0] r_V_149_reg_17211;
wire   [41:0] r_V_150_fu_531_p2;
reg   [41:0] r_V_150_reg_17215;
wire   [43:0] r_V_151_fu_517_p2;
reg   [43:0] r_V_151_reg_17219;
wire   [49:0] r_V_152_fu_516_p2;
reg   [49:0] r_V_152_reg_17223;
wire   [49:0] r_V_153_fu_473_p2;
reg   [49:0] r_V_153_reg_17227;
wire   [41:0] r_V_154_fu_523_p2;
reg   [41:0] r_V_154_reg_17231;
wire   [43:0] r_V_155_fu_483_p2;
reg   [43:0] r_V_155_reg_17235;
wire   [49:0] r_V_157_fu_467_p2;
reg   [49:0] r_V_157_reg_17239;
reg  signed [31:0] p_read_27_reg_41274;
reg  signed [31:0] p_read_27_reg_41274_pp0_iter1_reg;
reg  signed [31:0] p_read_27_reg_41274_pp0_iter2_reg;
reg  signed [31:0] p_read_28_reg_41284;
reg  signed [31:0] p_read_28_reg_41284_pp0_iter1_reg;
reg  signed [31:0] p_read_28_reg_41284_pp0_iter2_reg;
reg  signed [31:0] p_read_29_reg_41293;
reg  signed [31:0] p_read_29_reg_41293_pp0_iter1_reg;
reg  signed [31:0] p_read_30_reg_41303;
reg  signed [31:0] p_read_30_reg_41303_pp0_iter1_reg;
reg  signed [31:0] p_read_31_reg_41314;
reg  signed [31:0] p_read_32_reg_41324;
reg   [0:0] p_Result_s_reg_41333;
reg   [0:0] p_Result_403_reg_41339;
wire  signed [18:0] p_Val2_403_fu_17315_p2;
reg  signed [18:0] p_Val2_403_reg_41345;
reg   [0:0] p_Result_404_reg_41350;
reg   [0:0] Range2_all_ones_reg_41357;
reg   [0:0] p_Result_405_reg_41364;
reg   [0:0] p_Result_406_reg_41370;
wire  signed [19:0] p_Val2_406_fu_17379_p2;
reg  signed [19:0] p_Val2_406_reg_41376;
reg   [0:0] p_Result_407_reg_41381;
reg   [0:0] Range2_all_ones_79_reg_41388;
reg   [0:0] p_Result_408_reg_41395;
reg   [0:0] p_Result_409_reg_41401;
wire  signed [20:0] p_Val2_409_fu_17443_p2;
reg  signed [20:0] p_Val2_409_reg_41407;
reg   [0:0] p_Result_410_reg_41412;
reg   [0:0] Range2_all_ones_80_reg_41419;
reg   [0:0] p_Result_411_reg_41426;
reg   [0:0] p_Result_412_reg_41432;
wire  signed [18:0] p_Val2_412_fu_17507_p2;
reg  signed [18:0] p_Val2_412_reg_41438;
reg   [0:0] p_Result_413_reg_41443;
reg   [0:0] Range2_all_ones_81_reg_41450;
reg   [0:0] p_Result_414_reg_41457;
reg   [0:0] p_Result_415_reg_41463;
wire  signed [18:0] p_Val2_415_fu_17571_p2;
reg  signed [18:0] p_Val2_415_reg_41469;
reg   [0:0] p_Result_416_reg_41474;
reg   [0:0] Range2_all_ones_82_reg_41481;
reg   [0:0] p_Result_417_reg_41488;
reg   [0:0] p_Result_418_reg_41494;
wire  signed [20:0] p_Val2_418_fu_17635_p2;
reg  signed [20:0] p_Val2_418_reg_41500;
reg   [0:0] p_Result_419_reg_41505;
reg   [0:0] Range2_all_ones_83_reg_41512;
reg   [0:0] p_Result_420_reg_41519;
reg   [0:0] p_Result_421_reg_41525;
wire  signed [21:0] p_Val2_421_fu_17699_p2;
reg  signed [21:0] p_Val2_421_reg_41531;
reg   [0:0] p_Result_422_reg_41536;
reg   [0:0] Range2_all_ones_84_reg_41543;
reg   [0:0] p_Result_423_reg_41550;
reg   [0:0] p_Result_424_reg_41556;
wire  signed [16:0] p_Val2_424_fu_17763_p2;
reg  signed [16:0] p_Val2_424_reg_41562;
reg   [0:0] p_Result_425_reg_41567;
reg   [0:0] Range2_all_ones_85_reg_41574;
reg   [0:0] p_Result_426_reg_41581;
reg   [0:0] p_Result_427_reg_41587;
wire  signed [19:0] p_Val2_427_fu_17827_p2;
reg  signed [19:0] p_Val2_427_reg_41593;
reg   [0:0] p_Result_428_reg_41598;
reg   [0:0] Range2_all_ones_86_reg_41605;
reg   [0:0] p_Result_429_reg_41612;
reg   [20:0] p_Val2_429_reg_41618;
reg   [0:0] p_Result_430_reg_41623;
reg   [0:0] tmp_693_reg_41629;
reg   [0:0] Range2_all_ones_87_reg_41634;
reg   [0:0] p_Result_432_reg_41641;
reg   [17:0] p_Val2_432_reg_41647;
reg   [0:0] p_Result_433_reg_41652;
reg   [0:0] tmp_699_reg_41658;
reg   [0:0] Range2_all_ones_88_reg_41663;
reg   [0:0] p_Result_435_reg_41670;
reg   [15:0] p_Val2_435_reg_41676;
reg   [0:0] p_Result_436_reg_41681;
reg   [0:0] tmp_705_reg_41687;
reg   [0:0] Range2_all_ones_89_reg_41692;
reg   [0:0] p_Result_438_reg_41699;
reg   [19:0] p_Val2_438_reg_41705;
reg   [0:0] p_Result_439_reg_41710;
reg   [0:0] tmp_711_reg_41716;
reg   [0:0] Range2_all_ones_90_reg_41721;
reg   [0:0] p_Result_441_reg_41728;
reg   [17:0] p_Val2_441_reg_41734;
reg   [0:0] p_Result_442_reg_41739;
reg   [0:0] tmp_717_reg_41745;
reg   [0:0] Range2_all_ones_91_reg_41750;
wire  signed [16:0] p_Val2_445_fu_18169_p2;
reg  signed [16:0] p_Val2_445_reg_41757;
wire   [0:0] overflow_175_fu_18271_p2;
reg   [0:0] overflow_175_reg_41762;
wire   [0:0] or_ln346_94_fu_18301_p2;
reg   [0:0] or_ln346_94_reg_41767;
reg   [0:0] p_Result_447_reg_41772;
reg   [17:0] p_Val2_447_reg_41778;
reg   [0:0] p_Result_448_reg_41783;
reg   [0:0] tmp_729_reg_41789;
reg   [0:0] Range2_all_ones_93_reg_41794;
reg   [0:0] p_Result_450_reg_41801;
reg   [18:0] p_Val2_450_reg_41807;
reg   [0:0] p_Result_451_reg_41812;
reg   [0:0] tmp_735_reg_41818;
reg   [0:0] Range2_all_ones_94_reg_41823;
reg   [0:0] p_Result_453_reg_41830;
reg   [14:0] p_Val2_453_reg_41836;
reg   [0:0] p_Result_454_reg_41841;
reg   [0:0] tmp_741_reg_41847;
reg   [0:0] Range2_all_ones_95_reg_41852;
reg   [0:0] p_Result_456_reg_41859;
reg   [30:0] p_Val2_456_reg_41865;
reg   [0:0] p_Result_457_reg_41870;
reg   [0:0] tmp_747_reg_41876;
reg   [0:0] Range2_all_ones_96_reg_41881;
reg   [0:0] p_Result_459_reg_41888;
reg   [19:0] p_Val2_459_reg_41894;
reg   [0:0] p_Result_460_reg_41899;
reg   [0:0] tmp_753_reg_41905;
reg   [0:0] Range2_all_ones_97_reg_41910;
reg   [0:0] p_Result_462_reg_41917;
reg   [16:0] p_Val2_462_reg_41923;
reg   [0:0] p_Result_463_reg_41928;
reg   [0:0] tmp_759_reg_41934;
reg   [0:0] Range2_all_ones_98_reg_41939;
reg   [0:0] p_Result_465_reg_41946;
reg   [31:0] p_Val2_465_reg_41952;
reg   [0:0] p_Result_466_reg_41957;
reg   [0:0] tmp_765_reg_41963;
reg   [0:0] Range2_all_ones_99_reg_41968;
reg   [0:0] p_Result_468_reg_41975;
reg   [27:0] p_Val2_468_reg_41981;
reg   [0:0] p_Result_469_reg_41986;
reg   [0:0] tmp_771_reg_41992;
reg   [0:0] Range2_all_ones_100_reg_41997;
reg   [0:0] p_Result_471_reg_42004;
reg   [20:0] p_Val2_471_reg_42010;
reg   [0:0] p_Result_472_reg_42015;
reg   [0:0] tmp_777_reg_42021;
reg   [0:0] Range2_all_ones_101_reg_42026;
reg   [0:0] p_Result_474_reg_42033;
reg   [18:0] p_Val2_474_reg_42039;
reg   [0:0] p_Result_475_reg_42044;
reg   [0:0] tmp_783_reg_42050;
reg   [0:0] Range2_all_ones_102_reg_42055;
reg   [0:0] p_Result_477_reg_42062;
reg   [16:0] p_Val2_477_reg_42068;
reg   [0:0] p_Result_478_reg_42073;
reg   [0:0] tmp_789_reg_42079;
reg   [0:0] Range2_all_ones_103_reg_42084;
reg   [0:0] p_Result_480_reg_42091;
reg   [22:0] p_Val2_480_reg_42097;
reg   [0:0] p_Result_481_reg_42102;
reg   [0:0] tmp_795_reg_42108;
reg   [0:0] Range2_all_ones_104_reg_42113;
reg   [0:0] tmp_837_reg_42120;
reg   [0:0] tmp_909_reg_42125;
reg   [0:0] tmp_909_reg_42125_pp0_iter1_reg;
reg   [0:0] tmp_1011_reg_42130;
reg   [0:0] tmp_1011_reg_42130_pp0_iter1_reg;
wire  signed [31:0] rhs_98_fu_21437_p3;
reg  signed [31:0] rhs_98_reg_42135;
wire  signed [20:0] p_Val2_460_fu_21451_p2;
reg  signed [20:0] p_Val2_460_reg_42141;
wire   [0:0] overflow_180_fu_21539_p2;
reg   [0:0] overflow_180_reg_42146;
wire   [0:0] or_ln346_99_fu_21568_p2;
reg   [0:0] or_ln346_99_reg_42151;
wire  signed [17:0] p_Val2_463_fu_21580_p2;
reg  signed [17:0] p_Val2_463_reg_42156;
wire   [0:0] overflow_181_fu_21668_p2;
reg   [0:0] overflow_181_reg_42161;
wire   [0:0] or_ln346_100_fu_21697_p2;
reg   [0:0] or_ln346_100_reg_42166;
wire  signed [31:0] rhs_101_fu_21836_p3;
reg  signed [31:0] rhs_101_reg_42171;
wire  signed [28:0] p_Val2_469_fu_21850_p2;
reg  signed [28:0] p_Val2_469_reg_42177;
wire   [0:0] overflow_183_fu_21938_p2;
reg   [0:0] overflow_183_reg_42182;
wire   [0:0] or_ln346_102_fu_21967_p2;
reg   [0:0] or_ln346_102_reg_42187;
wire  signed [21:0] p_Val2_472_fu_21979_p2;
reg  signed [21:0] p_Val2_472_reg_42192;
wire   [0:0] overflow_184_fu_22067_p2;
reg   [0:0] overflow_184_reg_42197;
wire   [0:0] or_ln346_103_fu_22096_p2;
reg   [0:0] or_ln346_103_reg_42202;
wire  signed [19:0] p_Val2_475_fu_22108_p2;
reg  signed [19:0] p_Val2_475_reg_42207;
wire   [0:0] overflow_185_fu_22196_p2;
reg   [0:0] overflow_185_reg_42212;
wire   [0:0] or_ln346_104_fu_22225_p2;
reg   [0:0] or_ln346_104_reg_42217;
wire  signed [17:0] p_Val2_478_fu_22237_p2;
reg  signed [17:0] p_Val2_478_reg_42222;
wire   [0:0] overflow_186_fu_22325_p2;
reg   [0:0] overflow_186_reg_42227;
wire   [0:0] or_ln346_105_fu_22354_p2;
reg   [0:0] or_ln346_105_reg_42232;
wire  signed [23:0] p_Val2_481_fu_22366_p2;
reg  signed [23:0] p_Val2_481_reg_42237;
wire   [0:0] overflow_187_fu_22454_p2;
reg   [0:0] overflow_187_reg_42242;
wire   [0:0] or_ln346_106_fu_22483_p2;
reg   [0:0] or_ln346_106_reg_42247;
reg   [0:0] p_Result_483_reg_42252;
reg   [0:0] p_Result_484_reg_42258;
wire  signed [18:0] p_Val2_484_fu_22548_p2;
reg  signed [18:0] p_Val2_484_reg_42264;
reg   [0:0] p_Result_485_reg_42269;
reg   [0:0] Range2_all_ones_105_reg_42276;
reg   [0:0] p_Result_486_reg_42283;
reg   [0:0] p_Result_487_reg_42289;
wire  signed [19:0] p_Val2_487_fu_22612_p2;
reg  signed [19:0] p_Val2_487_reg_42295;
reg   [0:0] p_Result_488_reg_42300;
reg   [0:0] Range2_all_ones_106_reg_42307;
reg   [0:0] p_Result_489_reg_42314;
reg   [0:0] p_Result_490_reg_42320;
wire  signed [18:0] p_Val2_490_fu_22676_p2;
reg  signed [18:0] p_Val2_490_reg_42326;
reg   [0:0] p_Result_491_reg_42331;
reg   [0:0] Range2_all_ones_107_reg_42338;
reg   [0:0] p_Result_492_reg_42345;
reg   [0:0] p_Result_493_reg_42351;
wire  signed [19:0] p_Val2_493_fu_22740_p2;
reg  signed [19:0] p_Val2_493_reg_42357;
reg   [0:0] p_Result_494_reg_42362;
reg   [0:0] Range2_all_ones_108_reg_42369;
reg   [0:0] p_Result_495_reg_42376;
reg   [0:0] p_Result_496_reg_42382;
wire  signed [20:0] p_Val2_496_fu_22804_p2;
reg  signed [20:0] p_Val2_496_reg_42388;
reg   [0:0] p_Result_497_reg_42393;
reg   [0:0] Range2_all_ones_109_reg_42400;
reg   [0:0] p_Result_498_reg_42407;
reg   [0:0] p_Result_499_reg_42413;
wire  signed [18:0] p_Val2_499_fu_22868_p2;
reg  signed [18:0] p_Val2_499_reg_42419;
reg   [0:0] p_Result_500_reg_42424;
reg   [0:0] Range2_all_ones_110_reg_42431;
wire  signed [15:0] p_Val2_502_fu_22951_p2;
reg  signed [15:0] p_Val2_502_reg_42438;
wire   [0:0] overflow_194_fu_23053_p2;
reg   [0:0] overflow_194_reg_42443;
wire   [0:0] or_ln346_113_fu_23083_p2;
reg   [0:0] or_ln346_113_reg_42448;
reg   [0:0] p_Result_504_reg_42453;
reg   [0:0] p_Result_505_reg_42459;
wire  signed [20:0] p_Val2_505_fu_23131_p2;
reg  signed [20:0] p_Val2_505_reg_42465;
reg   [0:0] p_Result_506_reg_42470;
reg   [0:0] Range2_all_ones_112_reg_42477;
reg   [0:0] p_Result_507_reg_42484;
reg   [0:0] p_Result_508_reg_42490;
wire  signed [19:0] p_Val2_508_fu_23195_p2;
reg  signed [19:0] p_Val2_508_reg_42496;
reg   [0:0] p_Result_509_reg_42501;
reg   [0:0] Range2_all_ones_113_reg_42508;
reg   [0:0] p_Result_510_reg_42515;
reg   [30:0] p_Val2_510_reg_42521;
reg   [0:0] p_Result_511_reg_42526;
reg   [0:0] tmp_855_reg_42532;
reg   [0:0] Range2_all_ones_114_reg_42537;
reg   [0:0] p_Result_513_reg_42544;
reg   [17:0] p_Val2_513_reg_42550;
reg   [0:0] p_Result_514_reg_42555;
reg   [0:0] tmp_861_reg_42561;
reg   [0:0] Range2_all_ones_115_reg_42566;
reg   [0:0] p_Result_516_reg_42573;
reg   [20:0] p_Val2_516_reg_42579;
reg   [0:0] p_Result_517_reg_42584;
reg   [0:0] tmp_867_reg_42590;
reg   [0:0] Range2_all_ones_116_reg_42595;
reg   [0:0] p_Result_519_reg_42602;
reg   [20:0] p_Val2_519_reg_42608;
reg   [0:0] p_Result_520_reg_42613;
reg   [0:0] tmp_873_reg_42619;
reg   [0:0] Range2_all_ones_117_reg_42624;
reg   [0:0] p_Result_522_reg_42631;
reg   [22:0] p_Val2_522_reg_42637;
reg   [0:0] p_Result_523_reg_42642;
reg   [0:0] tmp_879_reg_42648;
reg   [0:0] Range2_all_ones_118_reg_42653;
reg   [0:0] p_Result_525_reg_42660;
reg   [18:0] p_Val2_525_reg_42666;
reg   [0:0] p_Result_526_reg_42671;
reg   [0:0] tmp_885_reg_42677;
reg   [0:0] Range2_all_ones_119_reg_42682;
reg   [0:0] p_Result_528_reg_42689;
reg   [20:0] p_Val2_528_reg_42695;
reg   [0:0] p_Result_529_reg_42700;
reg   [0:0] tmp_891_reg_42706;
reg   [0:0] Range2_all_ones_120_reg_42711;
reg   [0:0] p_Result_531_reg_42718;
reg   [19:0] p_Val2_531_reg_42724;
reg   [0:0] p_Result_532_reg_42729;
reg   [0:0] tmp_897_reg_42735;
reg   [0:0] Range2_all_ones_121_reg_42740;
reg   [0:0] p_Result_534_reg_42747;
reg   [19:0] p_Val2_534_reg_42753;
reg   [0:0] p_Result_535_reg_42758;
reg   [0:0] tmp_903_reg_42764;
reg   [0:0] Range2_all_ones_122_reg_42769;
wire  signed [31:0] lhs_80_fu_24598_p3;
reg  signed [31:0] lhs_80_reg_42776;
wire  signed [31:0] lhs_81_fu_24700_p3;
reg  signed [31:0] lhs_81_reg_42782;
wire  signed [31:0] lhs_82_fu_24802_p3;
reg  signed [31:0] lhs_82_reg_42788;
wire  signed [31:0] lhs_83_fu_24904_p3;
reg  signed [31:0] lhs_83_reg_42794;
wire  signed [31:0] lhs_84_fu_25006_p3;
reg  signed [31:0] lhs_84_reg_42800;
wire  signed [31:0] lhs_85_fu_25108_p3;
reg  signed [31:0] lhs_85_reg_42806;
wire  signed [31:0] lhs_86_fu_25210_p3;
reg  signed [31:0] lhs_86_reg_42812;
wire  signed [31:0] lhs_87_fu_25312_p3;
reg  signed [31:0] lhs_87_reg_42818;
wire  signed [31:0] lhs_88_fu_25414_p3;
reg  signed [31:0] lhs_88_reg_42824;
wire  signed [17:0] p_Val2_538_fu_27979_p2;
reg  signed [17:0] p_Val2_538_reg_42830;
wire   [0:0] overflow_206_fu_28081_p2;
reg   [0:0] overflow_206_reg_42835;
wire   [0:0] or_ln346_125_fu_28111_p2;
reg   [0:0] or_ln346_125_reg_42840;
reg   [0:0] p_Result_540_reg_42845;
reg   [0:0] p_Result_541_reg_42851;
wire  signed [19:0] p_Val2_541_fu_28159_p2;
reg  signed [19:0] p_Val2_541_reg_42857;
reg   [0:0] p_Result_542_reg_42862;
reg   [0:0] Range2_all_ones_124_reg_42869;
reg   [0:0] p_Result_543_reg_42876;
reg   [0:0] p_Result_544_reg_42882;
wire  signed [20:0] p_Val2_544_fu_28223_p2;
reg  signed [20:0] p_Val2_544_reg_42888;
reg   [0:0] p_Result_545_reg_42893;
reg   [0:0] Range2_all_ones_125_reg_42900;
reg   [0:0] p_Result_546_reg_42907;
reg   [0:0] p_Result_547_reg_42913;
wire  signed [19:0] p_Val2_547_fu_28287_p2;
reg  signed [19:0] p_Val2_547_reg_42919;
reg   [0:0] p_Result_548_reg_42924;
reg   [0:0] Range2_all_ones_126_reg_42931;
reg   [0:0] p_Result_549_reg_42938;
reg   [0:0] p_Result_550_reg_42944;
wire  signed [20:0] p_Val2_550_fu_28351_p2;
reg  signed [20:0] p_Val2_550_reg_42950;
reg   [0:0] p_Result_551_reg_42955;
reg   [0:0] Range2_all_ones_127_reg_42962;
reg   [0:0] p_Result_552_reg_42969;
reg   [0:0] p_Result_553_reg_42975;
wire  signed [19:0] p_Val2_553_fu_28415_p2;
reg  signed [19:0] p_Val2_553_reg_42981;
reg   [0:0] p_Result_554_reg_42986;
reg   [0:0] Range2_all_ones_128_reg_42993;
reg   [0:0] p_Result_555_reg_43000;
reg   [0:0] p_Result_556_reg_43006;
wire  signed [21:0] p_Val2_556_fu_28479_p2;
reg  signed [21:0] p_Val2_556_reg_43012;
reg   [0:0] p_Result_557_reg_43017;
reg   [0:0] Range2_all_ones_129_reg_43024;
reg   [0:0] p_Result_558_reg_43031;
reg   [0:0] p_Result_559_reg_43037;
wire  signed [16:0] p_Val2_559_fu_28543_p2;
reg  signed [16:0] p_Val2_559_reg_43043;
reg   [0:0] p_Result_560_reg_43048;
reg   [0:0] Range2_all_ones_130_reg_43055;
reg   [0:0] p_Result_561_reg_43062;
reg   [0:0] p_Result_562_reg_43068;
wire  signed [18:0] p_Val2_562_fu_28607_p2;
reg  signed [18:0] p_Val2_562_reg_43074;
reg   [0:0] p_Result_563_reg_43079;
reg   [0:0] Range2_all_ones_131_reg_43086;
reg   [0:0] p_Result_564_reg_43093;
reg   [19:0] p_Val2_564_reg_43099;
reg   [0:0] p_Result_565_reg_43104;
reg   [0:0] tmp_963_reg_43110;
reg   [0:0] Range2_all_ones_132_reg_43115;
reg   [0:0] p_Result_567_reg_43122;
reg   [18:0] p_Val2_567_reg_43128;
reg   [0:0] p_Result_568_reg_43133;
reg   [0:0] tmp_969_reg_43139;
reg   [0:0] Range2_all_ones_133_reg_43144;
reg   [0:0] p_Result_570_reg_43151;
reg   [18:0] p_Val2_570_reg_43157;
reg   [0:0] p_Result_571_reg_43162;
reg   [0:0] tmp_975_reg_43168;
reg   [0:0] Range2_all_ones_134_reg_43173;
reg   [0:0] p_Result_573_reg_43180;
reg   [19:0] p_Val2_573_reg_43186;
reg   [0:0] p_Result_574_reg_43191;
reg   [0:0] tmp_981_reg_43197;
reg   [0:0] Range2_all_ones_135_reg_43202;
reg   [0:0] p_Result_576_reg_43209;
reg   [18:0] p_Val2_576_reg_43215;
reg   [0:0] p_Result_577_reg_43220;
reg   [0:0] tmp_987_reg_43226;
reg   [0:0] Range2_all_ones_136_reg_43231;
reg   [0:0] p_Result_579_reg_43238;
reg   [18:0] p_Val2_579_reg_43244;
reg   [0:0] p_Result_580_reg_43249;
reg   [0:0] tmp_993_reg_43255;
reg   [0:0] Range2_all_ones_137_reg_43260;
reg   [0:0] p_Result_582_reg_43267;
reg   [16:0] p_Val2_582_reg_43273;
reg   [0:0] p_Result_583_reg_43278;
reg   [0:0] tmp_999_reg_43284;
reg   [0:0] Range2_all_ones_138_reg_43289;
reg   [0:0] p_Result_585_reg_43296;
reg   [17:0] p_Val2_585_reg_43302;
reg   [0:0] p_Result_586_reg_43307;
reg   [0:0] tmp_1005_reg_43313;
reg   [0:0] Range2_all_ones_139_reg_43318;
wire  signed [17:0] p_Val2_589_fu_29046_p2;
reg  signed [17:0] p_Val2_589_reg_43325;
wire   [0:0] overflow_223_fu_29148_p2;
reg   [0:0] overflow_223_reg_43330;
wire   [0:0] or_ln346_142_fu_29178_p2;
reg   [0:0] or_ln346_142_reg_43335;
reg   [0:0] p_Result_717_reg_43340;
wire   [31:0] p_Val2_717_fu_31020_p2;
reg   [31:0] p_Val2_717_reg_43347;
reg   [0:0] p_Result_718_reg_43353;
reg   [0:0] p_Result_719_reg_43360;
wire   [31:0] p_Val2_719_fu_31056_p2;
reg   [31:0] p_Val2_719_reg_43367;
reg   [0:0] p_Result_720_reg_43373;
reg   [0:0] p_Result_721_reg_43380;
wire   [31:0] p_Val2_721_fu_31092_p2;
reg   [31:0] p_Val2_721_reg_43387;
reg   [0:0] p_Result_722_reg_43393;
reg   [0:0] p_Result_723_reg_43400;
wire   [31:0] p_Val2_723_fu_31128_p2;
reg   [31:0] p_Val2_723_reg_43407;
reg   [0:0] p_Result_724_reg_43413;
reg   [0:0] p_Result_725_reg_43420;
wire   [31:0] p_Val2_725_fu_31164_p2;
reg   [31:0] p_Val2_725_reg_43427;
reg   [0:0] p_Result_726_reg_43433;
reg   [0:0] p_Result_727_reg_43440;
wire   [31:0] p_Val2_727_fu_31200_p2;
reg   [31:0] p_Val2_727_reg_43447;
reg   [0:0] p_Result_728_reg_43453;
reg   [0:0] p_Result_729_reg_43460;
wire   [31:0] p_Val2_729_fu_31236_p2;
reg   [31:0] p_Val2_729_reg_43467;
reg   [0:0] p_Result_730_reg_43473;
reg   [0:0] p_Result_731_reg_43480;
wire   [31:0] p_Val2_731_fu_31272_p2;
reg   [31:0] p_Val2_731_reg_43487;
reg   [0:0] p_Result_732_reg_43493;
reg   [0:0] p_Result_733_reg_43500;
wire   [31:0] p_Val2_733_fu_31308_p2;
reg   [31:0] p_Val2_733_reg_43507;
reg   [0:0] p_Result_734_reg_43513;
reg   [0:0] p_Result_591_reg_43520;
reg   [0:0] p_Result_592_reg_43526;
wire   [31:0] p_Val2_592_fu_33614_p2;
reg   [31:0] p_Val2_592_reg_43532;
reg   [0:0] p_Result_593_reg_43537;
reg   [0:0] Range2_all_ones_141_reg_43544;
reg   [0:0] p_Result_594_reg_43551;
reg   [0:0] p_Result_595_reg_43557;
wire  signed [20:0] p_Val2_595_fu_33678_p2;
reg  signed [20:0] p_Val2_595_reg_43563;
reg   [0:0] p_Result_596_reg_43568;
reg   [0:0] Range2_all_ones_142_reg_43575;
reg   [0:0] p_Result_597_reg_43582;
reg   [0:0] p_Result_598_reg_43588;
wire  signed [19:0] p_Val2_598_fu_33742_p2;
reg  signed [19:0] p_Val2_598_reg_43594;
reg   [0:0] p_Result_599_reg_43599;
reg   [0:0] Range2_all_ones_143_reg_43606;
reg   [0:0] p_Result_600_reg_43613;
reg   [0:0] p_Result_601_reg_43619;
wire  signed [26:0] p_Val2_601_fu_33806_p2;
reg  signed [26:0] p_Val2_601_reg_43625;
reg   [0:0] p_Result_602_reg_43630;
reg   [0:0] Range2_all_ones_144_reg_43637;
reg   [0:0] p_Result_603_reg_43644;
reg   [0:0] p_Result_604_reg_43650;
wire  signed [25:0] p_Val2_604_fu_33870_p2;
reg  signed [25:0] p_Val2_604_reg_43656;
reg   [0:0] p_Result_605_reg_43661;
reg   [0:0] Range2_all_ones_145_reg_43668;
reg   [0:0] p_Result_606_reg_43675;
reg   [0:0] p_Result_607_reg_43681;
wire  signed [20:0] p_Val2_607_fu_33934_p2;
reg  signed [20:0] p_Val2_607_reg_43687;
reg   [0:0] p_Result_608_reg_43692;
reg   [0:0] Range2_all_ones_146_reg_43699;
reg   [0:0] p_Result_609_reg_43706;
reg   [0:0] p_Result_610_reg_43712;
wire  signed [20:0] p_Val2_610_fu_33998_p2;
reg  signed [20:0] p_Val2_610_reg_43718;
reg   [0:0] p_Result_611_reg_43723;
reg   [0:0] Range2_all_ones_147_reg_43730;
reg   [0:0] p_Result_612_reg_43737;
reg   [0:0] p_Result_613_reg_43743;
wire  signed [20:0] p_Val2_613_fu_34062_p2;
reg  signed [20:0] p_Val2_613_reg_43749;
reg   [0:0] p_Result_614_reg_43754;
reg   [0:0] Range2_all_ones_148_reg_43761;
reg   [0:0] p_Result_615_reg_43768;
reg   [0:0] p_Result_616_reg_43774;
wire  signed [25:0] p_Val2_616_fu_34126_p2;
reg  signed [25:0] p_Val2_616_reg_43780;
reg   [0:0] p_Result_617_reg_43785;
reg   [0:0] Range2_all_ones_149_reg_43792;
reg   [0:0] p_Result_618_reg_43799;
reg   [30:0] p_Val2_618_reg_43805;
reg   [0:0] p_Result_619_reg_43810;
reg   [0:0] tmp_1071_reg_43816;
reg   [0:0] Range2_all_ones_150_reg_43821;
reg   [0:0] p_Result_621_reg_43828;
reg   [17:0] p_Val2_621_reg_43834;
reg   [0:0] p_Result_622_reg_43839;
reg   [0:0] tmp_1077_reg_43845;
reg   [0:0] Range2_all_ones_151_reg_43850;
reg   [0:0] p_Result_624_reg_43857;
reg   [19:0] p_Val2_624_reg_43863;
reg   [0:0] p_Result_625_reg_43868;
reg   [0:0] tmp_1083_reg_43874;
reg   [0:0] Range2_all_ones_152_reg_43879;
reg   [0:0] p_Result_627_reg_43886;
reg   [25:0] p_Val2_627_reg_43892;
reg   [0:0] p_Result_628_reg_43897;
reg   [0:0] tmp_1089_reg_43903;
reg   [0:0] Range2_all_ones_153_reg_43908;
reg   [0:0] p_Result_630_reg_43915;
reg   [25:0] p_Val2_630_reg_43921;
reg   [0:0] p_Result_631_reg_43926;
reg   [0:0] tmp_1095_reg_43932;
reg   [0:0] Range2_all_ones_154_reg_43937;
reg   [0:0] p_Result_633_reg_43944;
reg   [17:0] p_Val2_633_reg_43950;
reg   [0:0] p_Result_634_reg_43955;
reg   [0:0] tmp_1101_reg_43961;
reg   [0:0] Range2_all_ones_155_reg_43966;
reg   [0:0] p_Result_636_reg_43973;
reg   [19:0] p_Val2_636_reg_43979;
reg   [0:0] p_Result_637_reg_43984;
reg   [0:0] tmp_1107_reg_43990;
reg   [0:0] Range2_all_ones_156_reg_43995;
wire  signed [12:0] p_Val2_640_fu_34538_p2;
reg  signed [12:0] p_Val2_640_reg_44002;
wire   [0:0] overflow_240_fu_34640_p2;
reg   [0:0] overflow_240_reg_44007;
wire   [0:0] or_ln346_159_fu_34670_p2;
reg   [0:0] or_ln346_159_reg_44012;
reg   [0:0] p_Result_642_reg_44017;
reg   [25:0] p_Val2_642_reg_44023;
reg   [0:0] p_Result_643_reg_44028;
reg   [0:0] tmp_1119_reg_44034;
reg   [0:0] Range2_all_ones_158_reg_44039;
wire  signed [31:0] lhs_125_fu_36252_p3;
reg  signed [31:0] lhs_125_reg_44046;
wire  signed [31:0] lhs_126_fu_36354_p3;
reg  signed [31:0] lhs_126_reg_44052;
wire  signed [31:0] lhs_127_fu_36456_p3;
reg  signed [31:0] lhs_127_reg_44058;
wire  signed [31:0] lhs_128_fu_36558_p3;
reg  signed [31:0] lhs_128_reg_44064;
wire  signed [31:0] lhs_129_fu_36660_p3;
reg  signed [31:0] lhs_129_reg_44070;
wire  signed [31:0] lhs_130_fu_36762_p3;
reg  signed [31:0] lhs_130_reg_44076;
wire  signed [31:0] lhs_131_fu_36864_p3;
reg  signed [31:0] lhs_131_reg_44082;
wire  signed [31:0] lhs_132_fu_36966_p3;
reg  signed [31:0] lhs_132_reg_44088;
wire  signed [31:0] lhs_133_fu_37068_p3;
reg  signed [31:0] lhs_133_reg_44094;
wire  signed [31:0] r_V_124_fu_462_p0;
wire  signed [43:0] sext_ln70_74_fu_27903_p1;
wire   [11:0] r_V_124_fu_462_p1;
wire    ap_block_pp0_stage0;
wire  signed [31:0] r_V_107_fu_463_p0;
wire  signed [42:0] sext_ln70_64_fu_22494_p1;
wire  signed [10:0] r_V_107_fu_463_p1;
wire  signed [8:0] r_V_137_fu_464_p1;
wire  signed [20:0] r_V_99_fu_465_p1;
wire  signed [31:0] r_V_104_fu_466_p0;
wire  signed [41:0] sext_ln70_65_fu_22500_p1;
wire  signed [9:0] r_V_104_fu_466_p1;
wire  signed [31:0] r_V_157_fu_467_p0;
wire  signed [49:0] sext_ln70_86_fu_34148_p1;
wire  signed [17:0] r_V_157_fu_467_p1;
wire  signed [31:0] r_V_115_fu_468_p0;
wire  signed [44:0] sext_ln70_69_fu_23230_p1;
wire  signed [12:0] r_V_115_fu_468_p1;
wire  signed [14:0] r_V_103_fu_469_p1;
wire  signed [10:0] r_V_118_fu_470_p1;
wire  signed [31:0] r_V_112_fu_471_p0;
wire   [10:0] r_V_112_fu_471_p1;
wire  signed [31:0] r_V_123_fu_472_p0;
wire  signed [42:0] sext_ln70_75_fu_27908_p1;
wire   [10:0] r_V_123_fu_472_p1;
wire  signed [31:0] r_V_153_fu_473_p0;
wire  signed [17:0] r_V_153_fu_473_p1;
wire  signed [31:0] r_V_102_fu_474_p0;
wire  signed [40:0] sext_ln70_60_fu_18458_p1;
wire   [8:0] r_V_102_fu_474_p1;
wire  signed [9:0] r_V_114_fu_475_p1;
wire  signed [31:0] r_V_145_fu_476_p0;
wire  signed [43:0] sext_ln70_84_fu_33561_p1;
wire  signed [11:0] r_V_145_fu_476_p1;
wire  signed [31:0] r_V_121_fu_477_p0;
wire  signed [43:0] sext_ln70_66_fu_23217_p1;
wire  signed [11:0] r_V_121_fu_477_p1;
wire   [10:0] r_V_101_fu_478_p1;
wire  signed [31:0] r_V_127_fu_479_p0;
wire   [10:0] r_V_127_fu_479_p1;
wire  signed [31:0] r_V_90_fu_480_p0;
wire  signed [41:0] sext_ln70_53_fu_17869_p1;
wire  signed [9:0] r_V_90_fu_480_p1;
wire  signed [23:0] r_V_140_fu_481_p1;
wire  signed [11:0] r_V_89_fu_482_p1;
wire  signed [31:0] r_V_155_fu_483_p0;
wire  signed [43:0] sext_ln70_87_fu_34154_p1;
wire  signed [11:0] r_V_155_fu_483_p1;
wire  signed [31:0] r_V_79_fu_484_p0;
wire  signed [43:0] sext_ln70_46_fu_17254_p1;
wire  signed [11:0] r_V_79_fu_484_p1;
wire  signed [31:0] r_V_109_fu_485_p0;
wire   [9:0] r_V_109_fu_485_p1;
wire  signed [31:0] r_V_133_fu_486_p0;
wire  signed [42:0] sext_ln70_79_fu_28637_p1;
wire   [10:0] r_V_133_fu_486_p1;
wire  signed [31:0] r_V_81_fu_489_p0;
wire  signed [41:0] sext_ln70_48_fu_17266_p1;
wire   [9:0] r_V_81_fu_489_p1;
wire  signed [31:0] r_V_144_fu_490_p0;
wire  signed [48:0] sext_ln70_81_fu_33548_p1;
wire   [16:0] r_V_144_fu_490_p1;
wire  signed [9:0] r_V_130_fu_491_p1;
wire  signed [10:0] r_V_142_fu_492_p1;
wire   [23:0] r_V_149_fu_493_p1;
wire  signed [7:0] r_V_84_fu_494_p1;
wire  signed [31:0] r_V_85_fu_495_p0;
wire  signed [42:0] sext_ln70_47_fu_17260_p1;
wire   [10:0] r_V_85_fu_495_p1;
wire  signed [31:0] r_V_135_fu_496_p0;
wire   [10:0] r_V_135_fu_496_p1;
wire  signed [31:0] r_V_82_fu_497_p0;
wire  signed [11:0] r_V_82_fu_497_p1;
wire  signed [7:0] r_V_88_fu_498_p1;
wire  signed [6:0] r_V_94_fu_499_p1;
wire  signed [31:0] r_V_136_fu_500_p0;
wire  signed [10:0] r_V_136_fu_500_p1;
wire   [24:0] r_V_98_fu_501_p1;
wire  signed [23:0] r_V_95_fu_503_p1;
wire  signed [31:0] r_V_97_fu_504_p0;
wire   [8:0] r_V_97_fu_504_p1;
wire   [12:0] r_V_86_fu_505_p1;
wire  signed [31:0] r_V_131_fu_506_p0;
wire  signed [43:0] sext_ln70_80_fu_28644_p1;
wire  signed [11:0] r_V_131_fu_506_p1;
wire   [12:0] r_V_83_fu_507_p1;
wire  signed [31:0] r_V_147_fu_508_p0;
wire   [11:0] r_V_147_fu_508_p1;
wire  signed [31:0] r_V_80_fu_509_p0;
wire   [9:0] r_V_80_fu_509_p1;
wire  signed [31:0] r_V_125_fu_510_p0;
wire   [10:0] r_V_125_fu_510_p1;
wire  signed [31:0] r_V_106_fu_512_p0;
wire  signed [9:0] r_V_106_fu_512_p1;
wire   [12:0] r_V_128_fu_513_p1;
wire  signed [31:0] r_V_146_fu_514_p0;
wire   [11:0] r_V_146_fu_514_p1;
wire  signed [31:0] r_V_126_fu_515_p0;
wire  signed [11:0] r_V_126_fu_515_p1;
wire  signed [31:0] r_V_152_fu_516_p0;
wire   [17:0] r_V_152_fu_516_p1;
wire  signed [31:0] r_V_151_fu_517_p0;
wire  signed [11:0] r_V_151_fu_517_p1;
wire  signed [31:0] r_V_148_fu_518_p0;
wire   [16:0] r_V_148_fu_518_p1;
wire  signed [14:0] r_V_117_fu_519_p1;
wire  signed [31:0] r_V_120_fu_520_p0;
wire   [11:0] r_V_120_fu_520_p1;
wire   [7:0] r_V_129_fu_521_p1;
wire  signed [31:0] r_V_92_fu_522_p0;
wire   [9:0] r_V_92_fu_522_p1;
wire  signed [31:0] r_V_154_fu_523_p0;
wire  signed [41:0] sext_ln70_88_fu_34159_p1;
wire   [9:0] r_V_154_fu_523_p1;
wire  signed [31:0] r_V_134_fu_525_p0;
wire  signed [11:0] r_V_134_fu_525_p1;
wire  signed [31:0] r_V_111_fu_526_p0;
wire  signed [43:0] sext_ln70_63_fu_22489_p1;
wire   [11:0] r_V_111_fu_526_p1;
wire  signed [31:0] r_V_78_fu_527_p0;
wire  signed [10:0] r_V_78_fu_527_p1;
wire   [9:0] r_V_138_fu_528_p1;
wire  signed [31:0] r_V_108_fu_529_p0;
wire   [11:0] r_V_108_fu_529_p1;
wire   [11:0] r_V_96_fu_530_p1;
wire  signed [31:0] r_V_150_fu_531_p0;
wire   [9:0] r_V_150_fu_531_p1;
wire   [10:0] r_V_93_fu_532_p1;
wire  signed [31:0] r_V_132_fu_533_p0;
wire  signed [10:0] r_V_132_fu_533_p1;
wire  signed [12:0] r_V_100_fu_534_p1;
wire   [23:0] r_V_113_fu_535_p1;
wire  signed [31:0] r_V_fu_536_p0;
wire   [9:0] r_V_fu_536_p1;
wire  signed [31:0] r_V_116_fu_537_p0;
wire  signed [12:0] r_V_116_fu_537_p1;
wire  signed [31:0] r_V_87_fu_538_p0;
wire   [9:0] r_V_87_fu_538_p1;
wire  signed [31:0] r_V_105_fu_539_p0;
wire  signed [10:0] r_V_105_fu_539_p1;
wire  signed [17:0] r_V_143_fu_540_p1;
wire  signed [31:0] r_V_141_fu_541_p0;
wire  signed [11:0] r_V_141_fu_541_p1;
wire  signed [31:0] r_V_119_fu_542_p0;
wire   [12:0] r_V_119_fu_542_p1;
wire  signed [31:0] sext_ln70_46_fu_17254_p0;
wire  signed [31:0] sext_ln70_47_fu_17260_p0;
wire  signed [31:0] sext_ln70_48_fu_17266_p0;
wire   [17:0] p_Val2_402_fu_17281_p4;
wire   [0:0] tmp_fu_17303_p3;
wire   [18:0] zext_ln377_fu_17311_p1;
wire  signed [18:0] sext_ln823_fu_17291_p1;
wire   [18:0] p_Val2_405_fu_17345_p4;
wire   [0:0] tmp_645_fu_17367_p3;
wire   [19:0] zext_ln377_81_fu_17375_p1;
wire  signed [19:0] sext_ln823_78_fu_17355_p1;
wire   [19:0] p_Val2_408_fu_17409_p4;
wire   [0:0] tmp_651_fu_17431_p3;
wire   [20:0] zext_ln377_82_fu_17439_p1;
wire  signed [20:0] sext_ln823_79_fu_17419_p1;
wire   [17:0] p_Val2_411_fu_17473_p4;
wire   [0:0] tmp_657_fu_17495_p3;
wire   [18:0] zext_ln377_83_fu_17503_p1;
wire  signed [18:0] sext_ln823_80_fu_17483_p1;
wire   [17:0] p_Val2_414_fu_17537_p4;
wire   [0:0] tmp_663_fu_17559_p3;
wire   [18:0] zext_ln377_84_fu_17567_p1;
wire  signed [18:0] sext_ln823_81_fu_17547_p1;
wire   [19:0] p_Val2_417_fu_17601_p4;
wire   [0:0] tmp_669_fu_17623_p3;
wire   [20:0] zext_ln377_85_fu_17631_p1;
wire  signed [20:0] sext_ln823_82_fu_17611_p1;
wire   [20:0] p_Val2_420_fu_17665_p4;
wire   [0:0] tmp_675_fu_17687_p3;
wire   [21:0] zext_ln377_86_fu_17695_p1;
wire  signed [21:0] sext_ln823_83_fu_17675_p1;
wire   [15:0] p_Val2_423_fu_17729_p4;
wire   [0:0] tmp_681_fu_17751_p3;
wire   [16:0] zext_ln377_87_fu_17759_p1;
wire  signed [16:0] sext_ln823_84_fu_17739_p1;
wire   [18:0] p_Val2_426_fu_17793_p4;
wire   [0:0] tmp_687_fu_17815_p3;
wire   [19:0] zext_ln377_88_fu_17823_p1;
wire  signed [19:0] sext_ln823_85_fu_17803_p1;
wire  signed [31:0] sext_ln70_53_fu_17869_p0;
wire  signed [31:0] shl_ln_fu_18091_p1;
wire   [38:0] shl_ln_fu_18091_p3;
wire  signed [39:0] sext_ln1273_fu_18099_p1;
wire  signed [31:0] shl_ln1273_s_fu_18109_p1;
wire   [32:0] shl_ln1273_s_fu_18109_p3;
wire   [39:0] sub_ln1273_fu_18103_p2;
wire  signed [39:0] sext_ln1273_13_fu_18117_p1;
wire   [39:0] r_V_91_fu_18121_p2;
wire   [15:0] p_Val2_444_fu_18135_p4;
wire   [0:0] tmp_723_fu_18157_p3;
wire   [16:0] zext_ln377_94_fu_18165_p1;
wire  signed [16:0] sext_ln823_91_fu_18145_p1;
wire   [0:0] p_Result_446_fu_18175_p3;
wire   [0:0] p_Result_445_fu_18149_p3;
wire   [0:0] xor_ln896_270_fu_18183_p2;
wire   [0:0] xor_ln888_186_fu_18203_p2;
wire   [0:0] Range2_all_ones_92_fu_18195_p3;
wire   [0:0] or_ln888_94_fu_18209_p2;
wire   [0:0] tmp_726_fu_18221_p3;
wire   [0:0] xor_ln890_92_fu_18229_p2;
wire   [0:0] or_ln890_94_fu_18235_p2;
wire   [0:0] carry_187_fu_18189_p2;
wire   [0:0] deleted_zeros_91_fu_18215_p2;
wire   [0:0] xor_ln895_270_fu_18253_p2;
wire   [0:0] p_Result_444_fu_18127_p3;
wire   [0:0] or_ln895_94_fu_18259_p2;
wire   [0:0] xor_ln895_271_fu_18265_p2;
wire   [0:0] deleted_ones_175_fu_18241_p2;
wire   [0:0] xor_ln896_271_fu_18277_p2;
wire   [0:0] and_ln891_94_fu_18247_p2;
wire   [0:0] or_ln896_94_fu_18283_p2;
wire   [0:0] xor_ln896_499_fu_18289_p2;
wire   [0:0] underflow_175_fu_18295_p2;
wire  signed [31:0] sext_ln70_60_fu_18458_p0;
wire  signed [31:0] trunc_ln1273_fu_18852_p0;
wire   [17:0] trunc_ln1273_fu_18852_p1;
wire  signed [31:0] trunc_ln1273_7_fu_18864_p0;
wire   [22:0] trunc_ln1273_7_fu_18864_p1;
wire   [23:0] trunc_ln1273_2_fu_18868_p3;
wire   [23:0] trunc_ln5_fu_18856_p3;
wire   [23:0] sub_ln823_fu_18876_p2;
wire  signed [31:0] trunc_ln1273_8_fu_18890_p0;
wire   [15:0] trunc_ln1273_8_fu_18890_p1;
wire  signed [31:0] trunc_ln1273_9_fu_18902_p0;
wire   [22:0] trunc_ln1273_9_fu_18902_p1;
wire   [23:0] trunc_ln1273_4_fu_18906_p3;
wire   [23:0] trunc_ln1273_3_fu_18894_p3;
wire   [23:0] sub_ln823_2_fu_18914_p2;
wire  signed [31:0] trunc_ln1273_10_fu_18928_p0;
wire   [15:0] trunc_ln1273_10_fu_18928_p1;
wire  signed [31:0] trunc_ln1273_11_fu_18940_p0;
wire   [18:0] trunc_ln1273_11_fu_18940_p1;
wire   [23:0] trunc_ln1273_6_fu_18944_p3;
wire   [23:0] trunc_ln1273_5_fu_18932_p3;
wire   [23:0] sub_ln823_3_fu_18952_p2;
wire   [0:0] xor_ln896_fu_18969_p2;
wire   [0:0] xor_ln888_fu_18979_p2;
wire   [0:0] or_ln888_fu_18984_p2;
wire   [0:0] tmp_642_fu_18994_p3;
wire   [0:0] xor_ln890_fu_19002_p2;
wire   [0:0] or_ln890_fu_19008_p2;
wire   [0:0] carry_159_fu_18974_p2;
wire   [0:0] deleted_zeros_fu_18989_p2;
wire   [0:0] xor_ln895_fu_19024_p2;
wire   [0:0] or_ln895_fu_19030_p2;
wire   [0:0] xor_ln895_243_fu_19035_p2;
wire   [0:0] deleted_ones_fu_19014_p2;
wire   [0:0] xor_ln896_243_fu_19046_p2;
wire   [0:0] and_ln891_fu_19019_p2;
wire   [0:0] or_ln896_fu_19052_p2;
wire   [0:0] xor_ln896_485_fu_19058_p2;
wire   [0:0] overflow_fu_19040_p2;
wire   [0:0] underflow_fu_19064_p2;
wire   [0:0] or_ln346_fu_19077_p2;
wire   [31:0] select_ln346_fu_19069_p3;
wire  signed [31:0] sext_ln856_fu_18966_p1;
wire   [0:0] xor_ln896_244_fu_19094_p2;
wire   [0:0] xor_ln888_160_fu_19104_p2;
wire   [0:0] or_ln888_81_fu_19109_p2;
wire   [0:0] tmp_648_fu_19119_p3;
wire   [0:0] xor_ln890_79_fu_19127_p2;
wire   [0:0] or_ln890_81_fu_19133_p2;
wire   [0:0] carry_161_fu_19099_p2;
wire   [0:0] deleted_zeros_78_fu_19114_p2;
wire   [0:0] xor_ln895_244_fu_19149_p2;
wire   [0:0] or_ln895_81_fu_19155_p2;
wire   [0:0] xor_ln895_245_fu_19160_p2;
wire   [0:0] deleted_ones_162_fu_19139_p2;
wire   [0:0] xor_ln896_245_fu_19171_p2;
wire   [0:0] and_ln891_81_fu_19144_p2;
wire   [0:0] or_ln896_81_fu_19177_p2;
wire   [0:0] xor_ln896_486_fu_19183_p2;
wire   [0:0] overflow_162_fu_19165_p2;
wire   [0:0] underflow_162_fu_19189_p2;
wire   [0:0] or_ln346_81_fu_19202_p2;
wire   [31:0] select_ln346_163_fu_19194_p3;
wire  signed [31:0] sext_ln856_78_fu_19091_p1;
wire   [0:0] xor_ln896_246_fu_19219_p2;
wire   [0:0] xor_ln888_162_fu_19229_p2;
wire   [0:0] or_ln888_82_fu_19234_p2;
wire   [0:0] tmp_654_fu_19244_p3;
wire   [0:0] xor_ln890_80_fu_19252_p2;
wire   [0:0] or_ln890_82_fu_19258_p2;
wire   [0:0] carry_163_fu_19224_p2;
wire   [0:0] deleted_zeros_79_fu_19239_p2;
wire   [0:0] xor_ln895_246_fu_19274_p2;
wire   [0:0] or_ln895_82_fu_19280_p2;
wire   [0:0] xor_ln895_247_fu_19285_p2;
wire   [0:0] deleted_ones_163_fu_19264_p2;
wire   [0:0] xor_ln896_247_fu_19296_p2;
wire   [0:0] and_ln891_82_fu_19269_p2;
wire   [0:0] or_ln896_82_fu_19302_p2;
wire   [0:0] xor_ln896_487_fu_19308_p2;
wire   [0:0] overflow_163_fu_19290_p2;
wire   [0:0] underflow_163_fu_19314_p2;
wire   [0:0] or_ln346_82_fu_19327_p2;
wire   [31:0] select_ln346_164_fu_19319_p3;
wire  signed [31:0] sext_ln856_79_fu_19216_p1;
wire   [0:0] xor_ln896_248_fu_19344_p2;
wire   [0:0] xor_ln888_164_fu_19354_p2;
wire   [0:0] or_ln888_83_fu_19359_p2;
wire   [0:0] tmp_660_fu_19369_p3;
wire   [0:0] xor_ln890_81_fu_19377_p2;
wire   [0:0] or_ln890_83_fu_19383_p2;
wire   [0:0] carry_165_fu_19349_p2;
wire   [0:0] deleted_zeros_80_fu_19364_p2;
wire   [0:0] xor_ln895_248_fu_19399_p2;
wire   [0:0] or_ln895_83_fu_19405_p2;
wire   [0:0] xor_ln895_249_fu_19410_p2;
wire   [0:0] deleted_ones_164_fu_19389_p2;
wire   [0:0] xor_ln896_249_fu_19421_p2;
wire   [0:0] and_ln891_83_fu_19394_p2;
wire   [0:0] or_ln896_83_fu_19427_p2;
wire   [0:0] xor_ln896_488_fu_19433_p2;
wire   [0:0] overflow_164_fu_19415_p2;
wire   [0:0] underflow_164_fu_19439_p2;
wire   [0:0] or_ln346_83_fu_19452_p2;
wire   [31:0] select_ln346_165_fu_19444_p3;
wire  signed [31:0] sext_ln856_80_fu_19341_p1;
wire   [0:0] xor_ln896_250_fu_19469_p2;
wire   [0:0] xor_ln888_166_fu_19479_p2;
wire   [0:0] or_ln888_84_fu_19484_p2;
wire   [0:0] tmp_666_fu_19494_p3;
wire   [0:0] xor_ln890_82_fu_19502_p2;
wire   [0:0] or_ln890_84_fu_19508_p2;
wire   [0:0] carry_167_fu_19474_p2;
wire   [0:0] deleted_zeros_81_fu_19489_p2;
wire   [0:0] xor_ln895_250_fu_19524_p2;
wire   [0:0] or_ln895_84_fu_19530_p2;
wire   [0:0] xor_ln895_251_fu_19535_p2;
wire   [0:0] deleted_ones_165_fu_19514_p2;
wire   [0:0] xor_ln896_251_fu_19546_p2;
wire   [0:0] and_ln891_84_fu_19519_p2;
wire   [0:0] or_ln896_84_fu_19552_p2;
wire   [0:0] xor_ln896_489_fu_19558_p2;
wire   [0:0] overflow_165_fu_19540_p2;
wire   [0:0] underflow_165_fu_19564_p2;
wire   [0:0] or_ln346_84_fu_19577_p2;
wire   [31:0] select_ln346_166_fu_19569_p3;
wire  signed [31:0] sext_ln856_81_fu_19466_p1;
wire   [0:0] xor_ln896_252_fu_19594_p2;
wire   [0:0] xor_ln888_168_fu_19604_p2;
wire   [0:0] or_ln888_85_fu_19609_p2;
wire   [0:0] tmp_672_fu_19619_p3;
wire   [0:0] xor_ln890_83_fu_19627_p2;
wire   [0:0] or_ln890_85_fu_19633_p2;
wire   [0:0] carry_169_fu_19599_p2;
wire   [0:0] deleted_zeros_82_fu_19614_p2;
wire   [0:0] xor_ln895_252_fu_19649_p2;
wire   [0:0] or_ln895_85_fu_19655_p2;
wire   [0:0] xor_ln895_253_fu_19660_p2;
wire   [0:0] deleted_ones_166_fu_19639_p2;
wire   [0:0] xor_ln896_253_fu_19671_p2;
wire   [0:0] and_ln891_85_fu_19644_p2;
wire   [0:0] or_ln896_85_fu_19677_p2;
wire   [0:0] xor_ln896_490_fu_19683_p2;
wire   [0:0] overflow_166_fu_19665_p2;
wire   [0:0] underflow_166_fu_19689_p2;
wire   [0:0] or_ln346_85_fu_19702_p2;
wire   [31:0] select_ln346_167_fu_19694_p3;
wire  signed [31:0] sext_ln856_82_fu_19591_p1;
wire   [0:0] xor_ln896_254_fu_19719_p2;
wire   [0:0] xor_ln888_170_fu_19729_p2;
wire   [0:0] or_ln888_86_fu_19734_p2;
wire   [0:0] tmp_678_fu_19744_p3;
wire   [0:0] xor_ln890_84_fu_19752_p2;
wire   [0:0] or_ln890_86_fu_19758_p2;
wire   [0:0] carry_171_fu_19724_p2;
wire   [0:0] deleted_zeros_83_fu_19739_p2;
wire   [0:0] xor_ln895_254_fu_19774_p2;
wire   [0:0] or_ln895_86_fu_19780_p2;
wire   [0:0] xor_ln895_255_fu_19785_p2;
wire   [0:0] deleted_ones_167_fu_19764_p2;
wire   [0:0] xor_ln896_255_fu_19796_p2;
wire   [0:0] and_ln891_86_fu_19769_p2;
wire   [0:0] or_ln896_86_fu_19802_p2;
wire   [0:0] xor_ln896_491_fu_19808_p2;
wire   [0:0] overflow_167_fu_19790_p2;
wire   [0:0] underflow_167_fu_19814_p2;
wire   [0:0] or_ln346_86_fu_19827_p2;
wire   [31:0] select_ln346_168_fu_19819_p3;
wire  signed [31:0] sext_ln856_83_fu_19716_p1;
wire   [0:0] xor_ln896_256_fu_19844_p2;
wire   [0:0] xor_ln888_172_fu_19854_p2;
wire   [0:0] or_ln888_87_fu_19859_p2;
wire   [0:0] tmp_684_fu_19869_p3;
wire   [0:0] xor_ln890_85_fu_19877_p2;
wire   [0:0] or_ln890_87_fu_19883_p2;
wire   [0:0] carry_173_fu_19849_p2;
wire   [0:0] deleted_zeros_84_fu_19864_p2;
wire   [0:0] xor_ln895_256_fu_19899_p2;
wire   [0:0] or_ln895_87_fu_19905_p2;
wire   [0:0] xor_ln895_257_fu_19910_p2;
wire   [0:0] deleted_ones_168_fu_19889_p2;
wire   [0:0] xor_ln896_257_fu_19921_p2;
wire   [0:0] and_ln891_87_fu_19894_p2;
wire   [0:0] or_ln896_87_fu_19927_p2;
wire   [0:0] xor_ln896_492_fu_19933_p2;
wire   [0:0] overflow_168_fu_19915_p2;
wire   [0:0] underflow_168_fu_19939_p2;
wire   [0:0] or_ln346_87_fu_19952_p2;
wire   [31:0] select_ln346_169_fu_19944_p3;
wire  signed [31:0] sext_ln856_84_fu_19841_p1;
wire   [0:0] xor_ln896_258_fu_19969_p2;
wire   [0:0] xor_ln888_174_fu_19979_p2;
wire   [0:0] or_ln888_88_fu_19984_p2;
wire   [0:0] tmp_690_fu_19994_p3;
wire   [0:0] xor_ln890_86_fu_20002_p2;
wire   [0:0] or_ln890_88_fu_20008_p2;
wire   [0:0] carry_175_fu_19974_p2;
wire   [0:0] deleted_zeros_85_fu_19989_p2;
wire   [0:0] xor_ln895_258_fu_20024_p2;
wire   [0:0] or_ln895_88_fu_20030_p2;
wire   [0:0] xor_ln895_259_fu_20035_p2;
wire   [0:0] deleted_ones_169_fu_20014_p2;
wire   [0:0] xor_ln896_259_fu_20046_p2;
wire   [0:0] and_ln891_88_fu_20019_p2;
wire   [0:0] or_ln896_88_fu_20052_p2;
wire   [0:0] xor_ln896_493_fu_20058_p2;
wire   [0:0] overflow_169_fu_20040_p2;
wire   [0:0] underflow_169_fu_20064_p2;
wire   [0:0] or_ln346_88_fu_20077_p2;
wire   [31:0] select_ln346_170_fu_20069_p3;
wire  signed [31:0] sext_ln856_85_fu_19966_p1;
wire   [21:0] zext_ln377_89_fu_20094_p1;
wire  signed [21:0] sext_ln823_86_fu_20091_p1;
wire  signed [21:0] p_Val2_430_fu_20097_p2;
wire   [0:0] p_Result_431_fu_20107_p3;
wire   [0:0] xor_ln896_260_fu_20115_p2;
wire   [0:0] xor_ln888_176_fu_20126_p2;
wire   [0:0] or_ln888_89_fu_20131_p2;
wire   [0:0] tmp_696_fu_20142_p3;
wire   [0:0] xor_ln890_87_fu_20150_p2;
wire   [0:0] or_ln890_89_fu_20156_p2;
wire   [0:0] carry_177_fu_20121_p2;
wire   [0:0] deleted_zeros_86_fu_20137_p2;
wire   [0:0] xor_ln895_260_fu_20172_p2;
wire   [0:0] or_ln895_89_fu_20178_p2;
wire   [0:0] xor_ln895_261_fu_20184_p2;
wire   [0:0] deleted_ones_170_fu_20162_p2;
wire   [0:0] xor_ln896_261_fu_20195_p2;
wire   [0:0] and_ln891_89_fu_20167_p2;
wire   [0:0] or_ln896_89_fu_20201_p2;
wire   [0:0] xor_ln896_494_fu_20207_p2;
wire   [0:0] overflow_170_fu_20189_p2;
wire   [0:0] underflow_170_fu_20213_p2;
wire   [0:0] or_ln346_89_fu_20226_p2;
wire   [31:0] select_ln346_171_fu_20218_p3;
wire  signed [31:0] sext_ln856_86_fu_20103_p1;
wire   [18:0] zext_ln377_90_fu_20243_p1;
wire  signed [18:0] sext_ln823_87_fu_20240_p1;
wire  signed [18:0] p_Val2_433_fu_20246_p2;
wire   [0:0] p_Result_434_fu_20256_p3;
wire   [0:0] xor_ln896_262_fu_20264_p2;
wire   [0:0] xor_ln888_178_fu_20275_p2;
wire   [0:0] or_ln888_90_fu_20280_p2;
wire   [0:0] tmp_702_fu_20291_p3;
wire   [0:0] xor_ln890_88_fu_20299_p2;
wire   [0:0] or_ln890_90_fu_20305_p2;
wire   [0:0] carry_179_fu_20270_p2;
wire   [0:0] deleted_zeros_87_fu_20286_p2;
wire   [0:0] xor_ln895_262_fu_20321_p2;
wire   [0:0] or_ln895_90_fu_20327_p2;
wire   [0:0] xor_ln895_263_fu_20333_p2;
wire   [0:0] deleted_ones_171_fu_20311_p2;
wire   [0:0] xor_ln896_263_fu_20344_p2;
wire   [0:0] and_ln891_90_fu_20316_p2;
wire   [0:0] or_ln896_90_fu_20350_p2;
wire   [0:0] xor_ln896_495_fu_20356_p2;
wire   [0:0] overflow_171_fu_20338_p2;
wire   [0:0] underflow_171_fu_20362_p2;
wire   [0:0] or_ln346_90_fu_20375_p2;
wire   [31:0] select_ln346_172_fu_20367_p3;
wire  signed [31:0] sext_ln856_87_fu_20252_p1;
wire   [16:0] zext_ln377_91_fu_20392_p1;
wire  signed [16:0] sext_ln823_88_fu_20389_p1;
wire  signed [16:0] p_Val2_436_fu_20395_p2;
wire   [0:0] p_Result_437_fu_20405_p3;
wire   [0:0] xor_ln896_264_fu_20413_p2;
wire   [0:0] xor_ln888_180_fu_20424_p2;
wire   [0:0] or_ln888_91_fu_20429_p2;
wire   [0:0] tmp_708_fu_20440_p3;
wire   [0:0] xor_ln890_89_fu_20448_p2;
wire   [0:0] or_ln890_91_fu_20454_p2;
wire   [0:0] carry_181_fu_20419_p2;
wire   [0:0] deleted_zeros_88_fu_20435_p2;
wire   [0:0] xor_ln895_264_fu_20470_p2;
wire   [0:0] or_ln895_91_fu_20476_p2;
wire   [0:0] xor_ln895_265_fu_20482_p2;
wire   [0:0] deleted_ones_172_fu_20460_p2;
wire   [0:0] xor_ln896_265_fu_20493_p2;
wire   [0:0] and_ln891_91_fu_20465_p2;
wire   [0:0] or_ln896_91_fu_20499_p2;
wire   [0:0] xor_ln896_496_fu_20505_p2;
wire   [0:0] overflow_172_fu_20487_p2;
wire   [0:0] underflow_172_fu_20511_p2;
wire   [0:0] or_ln346_91_fu_20524_p2;
wire   [31:0] select_ln346_173_fu_20516_p3;
wire  signed [31:0] sext_ln856_88_fu_20401_p1;
wire   [20:0] zext_ln377_92_fu_20541_p1;
wire  signed [20:0] sext_ln823_89_fu_20538_p1;
wire  signed [20:0] p_Val2_439_fu_20544_p2;
wire   [0:0] p_Result_440_fu_20554_p3;
wire   [0:0] xor_ln896_266_fu_20562_p2;
wire   [0:0] xor_ln888_182_fu_20573_p2;
wire   [0:0] or_ln888_92_fu_20578_p2;
wire   [0:0] tmp_714_fu_20589_p3;
wire   [0:0] xor_ln890_90_fu_20597_p2;
wire   [0:0] or_ln890_92_fu_20603_p2;
wire   [0:0] carry_183_fu_20568_p2;
wire   [0:0] deleted_zeros_89_fu_20584_p2;
wire   [0:0] xor_ln895_266_fu_20619_p2;
wire   [0:0] or_ln895_92_fu_20625_p2;
wire   [0:0] xor_ln895_267_fu_20631_p2;
wire   [0:0] deleted_ones_173_fu_20609_p2;
wire   [0:0] xor_ln896_267_fu_20642_p2;
wire   [0:0] and_ln891_92_fu_20614_p2;
wire   [0:0] or_ln896_92_fu_20648_p2;
wire   [0:0] xor_ln896_497_fu_20654_p2;
wire   [0:0] overflow_173_fu_20636_p2;
wire   [0:0] underflow_173_fu_20660_p2;
wire   [0:0] or_ln346_92_fu_20673_p2;
wire   [31:0] select_ln346_174_fu_20665_p3;
wire  signed [31:0] sext_ln856_89_fu_20550_p1;
wire   [18:0] zext_ln377_93_fu_20690_p1;
wire  signed [18:0] sext_ln823_90_fu_20687_p1;
wire  signed [18:0] p_Val2_442_fu_20693_p2;
wire   [0:0] p_Result_443_fu_20703_p3;
wire   [0:0] xor_ln896_268_fu_20711_p2;
wire   [0:0] xor_ln888_184_fu_20722_p2;
wire   [0:0] or_ln888_93_fu_20727_p2;
wire   [0:0] tmp_720_fu_20738_p3;
wire   [0:0] xor_ln890_91_fu_20746_p2;
wire   [0:0] or_ln890_93_fu_20752_p2;
wire   [0:0] carry_185_fu_20717_p2;
wire   [0:0] deleted_zeros_90_fu_20733_p2;
wire   [0:0] xor_ln895_268_fu_20768_p2;
wire   [0:0] or_ln895_93_fu_20774_p2;
wire   [0:0] xor_ln895_269_fu_20780_p2;
wire   [0:0] deleted_ones_174_fu_20758_p2;
wire   [0:0] xor_ln896_269_fu_20791_p2;
wire   [0:0] and_ln891_93_fu_20763_p2;
wire   [0:0] or_ln896_93_fu_20797_p2;
wire   [0:0] xor_ln896_498_fu_20803_p2;
wire   [0:0] overflow_174_fu_20785_p2;
wire   [0:0] underflow_174_fu_20809_p2;
wire   [0:0] or_ln346_93_fu_20822_p2;
wire   [31:0] select_ln346_175_fu_20814_p3;
wire  signed [31:0] sext_ln856_90_fu_20699_p1;
wire   [31:0] select_ln346_176_fu_20839_p3;
wire  signed [31:0] sext_ln856_91_fu_20836_p1;
wire   [18:0] zext_ln377_95_fu_20856_p1;
wire  signed [18:0] sext_ln823_92_fu_20853_p1;
wire  signed [18:0] p_Val2_448_fu_20859_p2;
wire   [0:0] p_Result_449_fu_20869_p3;
wire   [0:0] xor_ln896_272_fu_20877_p2;
wire   [0:0] xor_ln888_188_fu_20888_p2;
wire   [0:0] or_ln888_95_fu_20893_p2;
wire   [0:0] tmp_732_fu_20904_p3;
wire   [0:0] xor_ln890_93_fu_20912_p2;
wire   [0:0] or_ln890_95_fu_20918_p2;
wire   [0:0] carry_189_fu_20883_p2;
wire   [0:0] deleted_zeros_92_fu_20899_p2;
wire   [0:0] xor_ln895_272_fu_20934_p2;
wire   [0:0] or_ln895_95_fu_20940_p2;
wire   [0:0] xor_ln895_273_fu_20946_p2;
wire   [0:0] deleted_ones_176_fu_20924_p2;
wire   [0:0] xor_ln896_273_fu_20957_p2;
wire   [0:0] and_ln891_95_fu_20929_p2;
wire   [0:0] or_ln896_95_fu_20963_p2;
wire   [0:0] xor_ln896_500_fu_20969_p2;
wire   [0:0] overflow_176_fu_20951_p2;
wire   [0:0] underflow_176_fu_20975_p2;
wire   [0:0] or_ln346_95_fu_20988_p2;
wire   [31:0] select_ln346_177_fu_20980_p3;
wire  signed [31:0] sext_ln856_92_fu_20865_p1;
wire   [19:0] zext_ln377_96_fu_21005_p1;
wire  signed [19:0] sext_ln823_93_fu_21002_p1;
wire  signed [19:0] p_Val2_451_fu_21008_p2;
wire   [0:0] p_Result_452_fu_21018_p3;
wire   [0:0] xor_ln896_274_fu_21026_p2;
wire   [0:0] xor_ln888_190_fu_21037_p2;
wire   [0:0] or_ln888_96_fu_21042_p2;
wire   [0:0] tmp_738_fu_21053_p3;
wire   [0:0] xor_ln890_94_fu_21061_p2;
wire   [0:0] or_ln890_96_fu_21067_p2;
wire   [0:0] carry_191_fu_21032_p2;
wire   [0:0] deleted_zeros_93_fu_21048_p2;
wire   [0:0] xor_ln895_274_fu_21083_p2;
wire   [0:0] or_ln895_96_fu_21089_p2;
wire   [0:0] xor_ln895_275_fu_21095_p2;
wire   [0:0] deleted_ones_177_fu_21073_p2;
wire   [0:0] xor_ln896_275_fu_21106_p2;
wire   [0:0] and_ln891_96_fu_21078_p2;
wire   [0:0] or_ln896_96_fu_21112_p2;
wire   [0:0] xor_ln896_501_fu_21118_p2;
wire   [0:0] overflow_177_fu_21100_p2;
wire   [0:0] underflow_177_fu_21124_p2;
wire   [0:0] or_ln346_96_fu_21137_p2;
wire   [31:0] select_ln346_178_fu_21129_p3;
wire  signed [31:0] sext_ln856_93_fu_21014_p1;
wire   [15:0] zext_ln377_97_fu_21154_p1;
wire  signed [15:0] sext_ln823_94_fu_21151_p1;
wire  signed [15:0] p_Val2_454_fu_21157_p2;
wire   [0:0] p_Result_455_fu_21167_p3;
wire   [0:0] xor_ln896_276_fu_21175_p2;
wire   [0:0] xor_ln888_192_fu_21186_p2;
wire   [0:0] or_ln888_97_fu_21191_p2;
wire   [0:0] tmp_744_fu_21202_p3;
wire   [0:0] xor_ln890_95_fu_21210_p2;
wire   [0:0] or_ln890_97_fu_21216_p2;
wire   [0:0] carry_193_fu_21181_p2;
wire   [0:0] deleted_zeros_94_fu_21197_p2;
wire   [0:0] xor_ln895_276_fu_21232_p2;
wire   [0:0] or_ln895_97_fu_21238_p2;
wire   [0:0] xor_ln895_277_fu_21244_p2;
wire   [0:0] deleted_ones_178_fu_21222_p2;
wire   [0:0] xor_ln896_277_fu_21255_p2;
wire   [0:0] and_ln891_97_fu_21227_p2;
wire   [0:0] or_ln896_97_fu_21261_p2;
wire   [0:0] xor_ln896_502_fu_21267_p2;
wire   [0:0] overflow_178_fu_21249_p2;
wire   [0:0] underflow_178_fu_21273_p2;
wire   [0:0] or_ln346_97_fu_21286_p2;
wire   [31:0] select_ln346_179_fu_21278_p3;
wire  signed [31:0] sext_ln856_94_fu_21163_p1;
wire   [31:0] zext_ln377_98_fu_21303_p1;
wire  signed [31:0] sext_ln818_fu_21300_p1;
wire   [31:0] p_Val2_457_fu_21306_p2;
wire   [0:0] p_Result_458_fu_21312_p3;
wire   [0:0] xor_ln896_278_fu_21320_p2;
wire   [0:0] xor_ln888_194_fu_21331_p2;
wire   [0:0] or_ln888_98_fu_21336_p2;
wire   [0:0] tmp_750_fu_21347_p3;
wire   [0:0] xor_ln890_96_fu_21355_p2;
wire   [0:0] or_ln890_98_fu_21361_p2;
wire   [0:0] carry_195_fu_21326_p2;
wire   [0:0] deleted_zeros_95_fu_21342_p2;
wire   [0:0] xor_ln895_278_fu_21377_p2;
wire   [0:0] or_ln895_98_fu_21383_p2;
wire   [0:0] xor_ln895_279_fu_21389_p2;
wire   [0:0] deleted_ones_179_fu_21367_p2;
wire   [0:0] xor_ln896_279_fu_21400_p2;
wire   [0:0] and_ln891_98_fu_21372_p2;
wire   [0:0] or_ln896_98_fu_21406_p2;
wire   [0:0] xor_ln896_503_fu_21412_p2;
wire   [0:0] overflow_179_fu_21394_p2;
wire   [0:0] underflow_179_fu_21418_p2;
wire   [0:0] or_ln346_98_fu_21431_p2;
wire   [31:0] select_ln346_180_fu_21423_p3;
wire   [20:0] zext_ln377_99_fu_21448_p1;
wire  signed [20:0] sext_ln823_95_fu_21445_p1;
wire   [0:0] p_Result_461_fu_21457_p3;
wire   [0:0] xor_ln896_280_fu_21465_p2;
wire   [0:0] xor_ln888_196_fu_21476_p2;
wire   [0:0] or_ln888_99_fu_21481_p2;
wire   [0:0] tmp_756_fu_21492_p3;
wire   [0:0] xor_ln890_97_fu_21500_p2;
wire   [0:0] or_ln890_99_fu_21506_p2;
wire   [0:0] carry_197_fu_21471_p2;
wire   [0:0] deleted_zeros_96_fu_21487_p2;
wire   [0:0] xor_ln895_280_fu_21522_p2;
wire   [0:0] or_ln895_99_fu_21528_p2;
wire   [0:0] xor_ln895_281_fu_21534_p2;
wire   [0:0] deleted_ones_180_fu_21512_p2;
wire   [0:0] xor_ln896_281_fu_21545_p2;
wire   [0:0] and_ln891_99_fu_21517_p2;
wire   [0:0] or_ln896_99_fu_21551_p2;
wire   [0:0] xor_ln896_504_fu_21557_p2;
wire   [0:0] underflow_180_fu_21563_p2;
wire   [17:0] zext_ln377_100_fu_21577_p1;
wire  signed [17:0] sext_ln823_96_fu_21574_p1;
wire   [0:0] p_Result_464_fu_21586_p3;
wire   [0:0] xor_ln896_282_fu_21594_p2;
wire   [0:0] xor_ln888_198_fu_21605_p2;
wire   [0:0] or_ln888_100_fu_21610_p2;
wire   [0:0] tmp_762_fu_21621_p3;
wire   [0:0] xor_ln890_98_fu_21629_p2;
wire   [0:0] or_ln890_100_fu_21635_p2;
wire   [0:0] carry_199_fu_21600_p2;
wire   [0:0] deleted_zeros_97_fu_21616_p2;
wire   [0:0] xor_ln895_282_fu_21651_p2;
wire   [0:0] or_ln895_100_fu_21657_p2;
wire   [0:0] xor_ln895_283_fu_21663_p2;
wire   [0:0] deleted_ones_181_fu_21641_p2;
wire   [0:0] xor_ln896_283_fu_21674_p2;
wire   [0:0] and_ln891_100_fu_21646_p2;
wire   [0:0] or_ln896_100_fu_21680_p2;
wire   [0:0] xor_ln896_505_fu_21686_p2;
wire   [0:0] underflow_181_fu_21692_p2;
wire   [31:0] zext_ln377_101_fu_21703_p1;
wire   [31:0] p_Val2_466_fu_21706_p2;
wire   [0:0] p_Result_467_fu_21711_p3;
wire   [0:0] xor_ln896_284_fu_21719_p2;
wire   [0:0] xor_ln888_200_fu_21730_p2;
wire   [0:0] or_ln888_101_fu_21735_p2;
wire   [0:0] tmp_768_fu_21746_p3;
wire   [0:0] xor_ln890_99_fu_21754_p2;
wire   [0:0] or_ln890_101_fu_21760_p2;
wire   [0:0] carry_201_fu_21725_p2;
wire   [0:0] deleted_zeros_98_fu_21741_p2;
wire   [0:0] xor_ln895_284_fu_21776_p2;
wire   [0:0] or_ln895_101_fu_21782_p2;
wire   [0:0] xor_ln895_285_fu_21788_p2;
wire   [0:0] deleted_ones_182_fu_21766_p2;
wire   [0:0] xor_ln896_285_fu_21799_p2;
wire   [0:0] and_ln891_101_fu_21771_p2;
wire   [0:0] or_ln896_101_fu_21805_p2;
wire   [0:0] xor_ln896_506_fu_21811_p2;
wire   [0:0] overflow_182_fu_21793_p2;
wire   [0:0] underflow_182_fu_21817_p2;
wire   [0:0] or_ln346_101_fu_21830_p2;
wire   [31:0] select_ln346_183_fu_21822_p3;
wire   [28:0] zext_ln377_102_fu_21847_p1;
wire  signed [28:0] sext_ln823_97_fu_21844_p1;
wire   [0:0] p_Result_470_fu_21856_p3;
wire   [0:0] xor_ln896_286_fu_21864_p2;
wire   [0:0] xor_ln888_202_fu_21875_p2;
wire   [0:0] or_ln888_102_fu_21880_p2;
wire   [0:0] tmp_774_fu_21891_p3;
wire   [0:0] xor_ln890_100_fu_21899_p2;
wire   [0:0] or_ln890_102_fu_21905_p2;
wire   [0:0] carry_203_fu_21870_p2;
wire   [0:0] deleted_zeros_99_fu_21886_p2;
wire   [0:0] xor_ln895_286_fu_21921_p2;
wire   [0:0] or_ln895_102_fu_21927_p2;
wire   [0:0] xor_ln895_287_fu_21933_p2;
wire   [0:0] deleted_ones_183_fu_21911_p2;
wire   [0:0] xor_ln896_287_fu_21944_p2;
wire   [0:0] and_ln891_102_fu_21916_p2;
wire   [0:0] or_ln896_102_fu_21950_p2;
wire   [0:0] xor_ln896_507_fu_21956_p2;
wire   [0:0] underflow_183_fu_21962_p2;
wire   [21:0] zext_ln377_103_fu_21976_p1;
wire  signed [21:0] sext_ln823_98_fu_21973_p1;
wire   [0:0] p_Result_473_fu_21985_p3;
wire   [0:0] xor_ln896_288_fu_21993_p2;
wire   [0:0] xor_ln888_204_fu_22004_p2;
wire   [0:0] or_ln888_103_fu_22009_p2;
wire   [0:0] tmp_780_fu_22020_p3;
wire   [0:0] xor_ln890_101_fu_22028_p2;
wire   [0:0] or_ln890_103_fu_22034_p2;
wire   [0:0] carry_205_fu_21999_p2;
wire   [0:0] deleted_zeros_100_fu_22015_p2;
wire   [0:0] xor_ln895_288_fu_22050_p2;
wire   [0:0] or_ln895_103_fu_22056_p2;
wire   [0:0] xor_ln895_289_fu_22062_p2;
wire   [0:0] deleted_ones_184_fu_22040_p2;
wire   [0:0] xor_ln896_289_fu_22073_p2;
wire   [0:0] and_ln891_103_fu_22045_p2;
wire   [0:0] or_ln896_103_fu_22079_p2;
wire   [0:0] xor_ln896_508_fu_22085_p2;
wire   [0:0] underflow_184_fu_22091_p2;
wire   [19:0] zext_ln377_104_fu_22105_p1;
wire  signed [19:0] sext_ln823_99_fu_22102_p1;
wire   [0:0] p_Result_476_fu_22114_p3;
wire   [0:0] xor_ln896_290_fu_22122_p2;
wire   [0:0] xor_ln888_206_fu_22133_p2;
wire   [0:0] or_ln888_104_fu_22138_p2;
wire   [0:0] tmp_786_fu_22149_p3;
wire   [0:0] xor_ln890_102_fu_22157_p2;
wire   [0:0] or_ln890_104_fu_22163_p2;
wire   [0:0] carry_207_fu_22128_p2;
wire   [0:0] deleted_zeros_101_fu_22144_p2;
wire   [0:0] xor_ln895_290_fu_22179_p2;
wire   [0:0] or_ln895_104_fu_22185_p2;
wire   [0:0] xor_ln895_291_fu_22191_p2;
wire   [0:0] deleted_ones_185_fu_22169_p2;
wire   [0:0] xor_ln896_291_fu_22202_p2;
wire   [0:0] and_ln891_104_fu_22174_p2;
wire   [0:0] or_ln896_104_fu_22208_p2;
wire   [0:0] xor_ln896_509_fu_22214_p2;
wire   [0:0] underflow_185_fu_22220_p2;
wire   [17:0] zext_ln377_105_fu_22234_p1;
wire  signed [17:0] sext_ln823_100_fu_22231_p1;
wire   [0:0] p_Result_479_fu_22243_p3;
wire   [0:0] xor_ln896_292_fu_22251_p2;
wire   [0:0] xor_ln888_208_fu_22262_p2;
wire   [0:0] or_ln888_105_fu_22267_p2;
wire   [0:0] tmp_792_fu_22278_p3;
wire   [0:0] xor_ln890_103_fu_22286_p2;
wire   [0:0] or_ln890_105_fu_22292_p2;
wire   [0:0] carry_209_fu_22257_p2;
wire   [0:0] deleted_zeros_102_fu_22273_p2;
wire   [0:0] xor_ln895_292_fu_22308_p2;
wire   [0:0] or_ln895_105_fu_22314_p2;
wire   [0:0] xor_ln895_293_fu_22320_p2;
wire   [0:0] deleted_ones_186_fu_22298_p2;
wire   [0:0] xor_ln896_293_fu_22331_p2;
wire   [0:0] and_ln891_105_fu_22303_p2;
wire   [0:0] or_ln896_105_fu_22337_p2;
wire   [0:0] xor_ln896_510_fu_22343_p2;
wire   [0:0] underflow_186_fu_22349_p2;
wire   [23:0] zext_ln377_106_fu_22363_p1;
wire  signed [23:0] sext_ln823_101_fu_22360_p1;
wire   [0:0] p_Result_482_fu_22372_p3;
wire   [0:0] xor_ln896_294_fu_22380_p2;
wire   [0:0] xor_ln888_210_fu_22391_p2;
wire   [0:0] or_ln888_106_fu_22396_p2;
wire   [0:0] tmp_798_fu_22407_p3;
wire   [0:0] xor_ln890_104_fu_22415_p2;
wire   [0:0] or_ln890_106_fu_22421_p2;
wire   [0:0] carry_211_fu_22386_p2;
wire   [0:0] deleted_zeros_103_fu_22402_p2;
wire   [0:0] xor_ln895_294_fu_22437_p2;
wire   [0:0] or_ln895_106_fu_22443_p2;
wire   [0:0] xor_ln895_295_fu_22449_p2;
wire   [0:0] deleted_ones_187_fu_22427_p2;
wire   [0:0] xor_ln896_295_fu_22460_p2;
wire   [0:0] and_ln891_106_fu_22432_p2;
wire   [0:0] or_ln896_106_fu_22466_p2;
wire   [0:0] xor_ln896_511_fu_22472_p2;
wire   [0:0] underflow_187_fu_22478_p2;
wire   [17:0] p_Val2_483_fu_22514_p4;
wire   [0:0] tmp_801_fu_22536_p3;
wire   [18:0] zext_ln377_107_fu_22544_p1;
wire  signed [18:0] sext_ln823_102_fu_22524_p1;
wire   [18:0] p_Val2_486_fu_22578_p4;
wire   [0:0] tmp_807_fu_22600_p3;
wire   [19:0] zext_ln377_108_fu_22608_p1;
wire  signed [19:0] sext_ln823_103_fu_22588_p1;
wire   [17:0] p_Val2_489_fu_22642_p4;
wire   [0:0] tmp_813_fu_22664_p3;
wire   [18:0] zext_ln377_109_fu_22672_p1;
wire  signed [18:0] sext_ln823_104_fu_22652_p1;
wire   [18:0] p_Val2_492_fu_22706_p4;
wire   [0:0] tmp_819_fu_22728_p3;
wire   [19:0] zext_ln377_110_fu_22736_p1;
wire  signed [19:0] sext_ln823_105_fu_22716_p1;
wire   [19:0] p_Val2_495_fu_22770_p4;
wire   [0:0] tmp_825_fu_22792_p3;
wire   [20:0] zext_ln377_111_fu_22800_p1;
wire  signed [20:0] sext_ln823_106_fu_22780_p1;
wire   [17:0] p_Val2_498_fu_22834_p4;
wire   [0:0] tmp_831_fu_22856_p3;
wire   [18:0] zext_ln377_112_fu_22864_p1;
wire  signed [18:0] sext_ln823_107_fu_22844_p1;
wire   [37:0] shl_ln1273_12_fu_22890_p3;
wire   [32:0] shl_ln1273_13_fu_22901_p3;
wire  signed [38:0] sext_ln1273_15_fu_22908_p1;
wire  signed [38:0] sext_ln1273_14_fu_22897_p1;
wire   [38:0] r_V_110_fu_22912_p2;
wire   [14:0] p_Val2_501_fu_22926_p4;
wire   [15:0] zext_ln377_113_fu_22948_p1;
wire  signed [15:0] sext_ln823_108_fu_22936_p1;
wire   [0:0] p_Result_503_fu_22957_p3;
wire   [0:0] p_Result_502_fu_22940_p3;
wire   [0:0] xor_ln896_308_fu_22965_p2;
wire   [0:0] xor_ln888_224_fu_22985_p2;
wire   [0:0] Range2_all_ones_111_fu_22977_p3;
wire   [0:0] or_ln888_113_fu_22991_p2;
wire   [0:0] tmp_840_fu_23003_p3;
wire   [0:0] xor_ln890_111_fu_23011_p2;
wire   [0:0] or_ln890_113_fu_23017_p2;
wire   [0:0] carry_225_fu_22971_p2;
wire   [0:0] deleted_zeros_110_fu_22997_p2;
wire   [0:0] xor_ln895_308_fu_23035_p2;
wire   [0:0] p_Result_501_fu_22918_p3;
wire   [0:0] or_ln895_113_fu_23041_p2;
wire   [0:0] xor_ln895_309_fu_23047_p2;
wire   [0:0] deleted_ones_194_fu_23023_p2;
wire   [0:0] xor_ln896_309_fu_23059_p2;
wire   [0:0] and_ln891_113_fu_23029_p2;
wire   [0:0] or_ln896_113_fu_23065_p2;
wire   [0:0] xor_ln896_518_fu_23071_p2;
wire   [0:0] underflow_194_fu_23077_p2;
wire   [19:0] p_Val2_504_fu_23097_p4;
wire   [0:0] tmp_843_fu_23119_p3;
wire   [20:0] zext_ln377_114_fu_23127_p1;
wire  signed [20:0] sext_ln823_109_fu_23107_p1;
wire   [18:0] p_Val2_507_fu_23161_p4;
wire   [0:0] tmp_849_fu_23183_p3;
wire   [19:0] zext_ln377_115_fu_23191_p1;
wire  signed [19:0] sext_ln823_110_fu_23171_p1;
wire  signed [31:0] rhs_fu_19083_p3;
wire  signed [32:0] sext_ln813_fu_23622_p1;
wire   [32:0] ret_V_fu_23626_p2;
wire   [31:0] p_Val2_645_fu_23640_p2;
wire   [0:0] p_Result_645_fu_23632_p3;
wire   [0:0] p_Result_646_fu_23646_p3;
wire   [0:0] xor_ln895_404_fu_23654_p2;
wire   [0:0] xor_ln896_404_fu_23666_p2;
wire   [0:0] xor_ln302_fu_23678_p2;
wire   [0:0] overflow_242_fu_23660_p2;
wire   [0:0] xor_ln302_162_fu_23684_p2;
wire   [0:0] underflow_242_fu_23672_p2;
wire   [0:0] or_ln302_fu_23690_p2;
wire   [31:0] select_ln302_fu_23696_p3;
wire   [31:0] select_ln350_fu_23704_p3;
wire  signed [31:0] rhs_81_fu_19208_p3;
wire  signed [32:0] sext_ln813_153_fu_23720_p1;
wire   [32:0] ret_V_81_fu_23724_p2;
wire   [31:0] p_Val2_647_fu_23738_p2;
wire   [0:0] p_Result_647_fu_23730_p3;
wire   [0:0] p_Result_648_fu_23744_p3;
wire   [0:0] xor_ln895_405_fu_23752_p2;
wire   [0:0] xor_ln896_405_fu_23764_p2;
wire   [0:0] xor_ln302_163_fu_23776_p2;
wire   [0:0] overflow_243_fu_23758_p2;
wire   [0:0] xor_ln302_164_fu_23782_p2;
wire   [0:0] underflow_243_fu_23770_p2;
wire   [0:0] or_ln302_81_fu_23788_p2;
wire   [31:0] select_ln302_163_fu_23794_p3;
wire   [31:0] select_ln350_81_fu_23802_p3;
wire  signed [31:0] rhs_82_fu_19333_p3;
wire  signed [32:0] sext_ln813_154_fu_23818_p1;
wire   [32:0] ret_V_82_fu_23822_p2;
wire   [31:0] p_Val2_649_fu_23836_p2;
wire   [0:0] p_Result_649_fu_23828_p3;
wire   [0:0] p_Result_650_fu_23842_p3;
wire   [0:0] xor_ln895_406_fu_23850_p2;
wire   [0:0] xor_ln896_406_fu_23862_p2;
wire   [0:0] xor_ln302_165_fu_23874_p2;
wire   [0:0] overflow_244_fu_23856_p2;
wire   [0:0] xor_ln302_166_fu_23880_p2;
wire   [0:0] underflow_244_fu_23868_p2;
wire   [0:0] or_ln302_82_fu_23886_p2;
wire   [31:0] select_ln302_165_fu_23892_p3;
wire   [31:0] select_ln350_82_fu_23900_p3;
wire  signed [31:0] rhs_83_fu_19458_p3;
wire  signed [32:0] sext_ln813_155_fu_23916_p1;
wire   [32:0] ret_V_83_fu_23920_p2;
wire   [31:0] p_Val2_651_fu_23934_p2;
wire   [0:0] p_Result_651_fu_23926_p3;
wire   [0:0] p_Result_652_fu_23940_p3;
wire   [0:0] xor_ln895_407_fu_23948_p2;
wire   [0:0] xor_ln896_407_fu_23960_p2;
wire   [0:0] xor_ln302_167_fu_23972_p2;
wire   [0:0] overflow_245_fu_23954_p2;
wire   [0:0] xor_ln302_168_fu_23978_p2;
wire   [0:0] underflow_245_fu_23966_p2;
wire   [0:0] or_ln302_83_fu_23984_p2;
wire   [31:0] select_ln302_167_fu_23990_p3;
wire   [31:0] select_ln350_83_fu_23998_p3;
wire  signed [31:0] rhs_84_fu_19583_p3;
wire  signed [32:0] sext_ln813_156_fu_24014_p1;
wire   [32:0] ret_V_84_fu_24018_p2;
wire   [31:0] p_Val2_653_fu_24032_p2;
wire   [0:0] p_Result_653_fu_24024_p3;
wire   [0:0] p_Result_654_fu_24038_p3;
wire   [0:0] xor_ln895_408_fu_24046_p2;
wire   [0:0] xor_ln896_408_fu_24058_p2;
wire   [0:0] xor_ln302_169_fu_24070_p2;
wire   [0:0] overflow_246_fu_24052_p2;
wire   [0:0] xor_ln302_170_fu_24076_p2;
wire   [0:0] underflow_246_fu_24064_p2;
wire   [0:0] or_ln302_84_fu_24082_p2;
wire   [31:0] select_ln302_169_fu_24088_p3;
wire   [31:0] select_ln350_84_fu_24096_p3;
wire  signed [31:0] rhs_85_fu_19708_p3;
wire  signed [32:0] sext_ln813_157_fu_24112_p1;
wire   [32:0] ret_V_85_fu_24116_p2;
wire   [31:0] p_Val2_655_fu_24130_p2;
wire   [0:0] p_Result_655_fu_24122_p3;
wire   [0:0] p_Result_656_fu_24136_p3;
wire   [0:0] xor_ln895_409_fu_24144_p2;
wire   [0:0] xor_ln896_409_fu_24156_p2;
wire   [0:0] xor_ln302_171_fu_24168_p2;
wire   [0:0] overflow_247_fu_24150_p2;
wire   [0:0] xor_ln302_172_fu_24174_p2;
wire   [0:0] underflow_247_fu_24162_p2;
wire   [0:0] or_ln302_85_fu_24180_p2;
wire   [31:0] select_ln302_171_fu_24186_p3;
wire   [31:0] select_ln350_85_fu_24194_p3;
wire  signed [31:0] rhs_86_fu_19833_p3;
wire  signed [32:0] sext_ln813_158_fu_24210_p1;
wire   [32:0] ret_V_86_fu_24214_p2;
wire   [31:0] p_Val2_657_fu_24228_p2;
wire   [0:0] p_Result_657_fu_24220_p3;
wire   [0:0] p_Result_658_fu_24234_p3;
wire   [0:0] xor_ln895_410_fu_24242_p2;
wire   [0:0] xor_ln896_410_fu_24254_p2;
wire   [0:0] xor_ln302_173_fu_24266_p2;
wire   [0:0] overflow_248_fu_24248_p2;
wire   [0:0] xor_ln302_174_fu_24272_p2;
wire   [0:0] underflow_248_fu_24260_p2;
wire   [0:0] or_ln302_86_fu_24278_p2;
wire   [31:0] select_ln302_173_fu_24284_p3;
wire   [31:0] select_ln350_86_fu_24292_p3;
wire  signed [31:0] rhs_87_fu_19958_p3;
wire  signed [32:0] sext_ln813_159_fu_24308_p1;
wire   [32:0] ret_V_87_fu_24312_p2;
wire   [31:0] p_Val2_659_fu_24326_p2;
wire   [0:0] p_Result_659_fu_24318_p3;
wire   [0:0] p_Result_660_fu_24332_p3;
wire   [0:0] xor_ln895_411_fu_24340_p2;
wire   [0:0] xor_ln896_411_fu_24352_p2;
wire   [0:0] xor_ln302_175_fu_24364_p2;
wire   [0:0] overflow_249_fu_24346_p2;
wire   [0:0] xor_ln302_176_fu_24370_p2;
wire   [0:0] underflow_249_fu_24358_p2;
wire   [0:0] or_ln302_87_fu_24376_p2;
wire   [31:0] select_ln302_175_fu_24382_p3;
wire   [31:0] select_ln350_87_fu_24390_p3;
wire  signed [31:0] rhs_88_fu_20083_p3;
wire  signed [32:0] sext_ln813_160_fu_24406_p1;
wire   [32:0] ret_V_88_fu_24410_p2;
wire   [31:0] p_Val2_661_fu_24424_p2;
wire   [0:0] p_Result_661_fu_24416_p3;
wire   [0:0] p_Result_662_fu_24430_p3;
wire   [0:0] xor_ln895_412_fu_24438_p2;
wire   [0:0] xor_ln896_412_fu_24450_p2;
wire   [0:0] xor_ln302_177_fu_24462_p2;
wire   [0:0] overflow_250_fu_24444_p2;
wire   [0:0] xor_ln302_178_fu_24468_p2;
wire   [0:0] underflow_250_fu_24456_p2;
wire   [0:0] or_ln302_88_fu_24474_p2;
wire   [31:0] select_ln302_177_fu_24480_p3;
wire   [31:0] select_ln350_88_fu_24488_p3;
wire  signed [31:0] lhs_fu_23712_p3;
wire  signed [31:0] rhs_89_fu_20232_p3;
wire  signed [32:0] sext_ln813_162_fu_24508_p1;
wire  signed [32:0] sext_ln813_161_fu_24504_p1;
wire   [32:0] ret_V_89_fu_24512_p2;
wire   [31:0] p_Val2_663_fu_24526_p2;
wire   [0:0] p_Result_663_fu_24518_p3;
wire   [0:0] p_Result_664_fu_24532_p3;
wire   [0:0] xor_ln895_413_fu_24540_p2;
wire   [0:0] xor_ln896_413_fu_24552_p2;
wire   [0:0] xor_ln302_179_fu_24564_p2;
wire   [0:0] overflow_251_fu_24546_p2;
wire   [0:0] xor_ln302_180_fu_24570_p2;
wire   [0:0] underflow_251_fu_24558_p2;
wire   [0:0] or_ln302_89_fu_24576_p2;
wire   [31:0] select_ln302_179_fu_24582_p3;
wire   [31:0] select_ln350_89_fu_24590_p3;
wire  signed [31:0] lhs_72_fu_23810_p3;
wire  signed [31:0] rhs_90_fu_20381_p3;
wire  signed [32:0] sext_ln813_164_fu_24610_p1;
wire  signed [32:0] sext_ln813_163_fu_24606_p1;
wire   [32:0] ret_V_90_fu_24614_p2;
wire   [31:0] p_Val2_665_fu_24628_p2;
wire   [0:0] p_Result_665_fu_24620_p3;
wire   [0:0] p_Result_666_fu_24634_p3;
wire   [0:0] xor_ln895_414_fu_24642_p2;
wire   [0:0] xor_ln896_414_fu_24654_p2;
wire   [0:0] xor_ln302_181_fu_24666_p2;
wire   [0:0] overflow_252_fu_24648_p2;
wire   [0:0] xor_ln302_182_fu_24672_p2;
wire   [0:0] underflow_252_fu_24660_p2;
wire   [0:0] or_ln302_90_fu_24678_p2;
wire   [31:0] select_ln302_181_fu_24684_p3;
wire   [31:0] select_ln350_90_fu_24692_p3;
wire  signed [31:0] lhs_73_fu_23908_p3;
wire  signed [31:0] rhs_91_fu_20530_p3;
wire  signed [32:0] sext_ln813_166_fu_24712_p1;
wire  signed [32:0] sext_ln813_165_fu_24708_p1;
wire   [32:0] ret_V_91_fu_24716_p2;
wire   [31:0] p_Val2_667_fu_24730_p2;
wire   [0:0] p_Result_667_fu_24722_p3;
wire   [0:0] p_Result_668_fu_24736_p3;
wire   [0:0] xor_ln895_415_fu_24744_p2;
wire   [0:0] xor_ln896_415_fu_24756_p2;
wire   [0:0] xor_ln302_183_fu_24768_p2;
wire   [0:0] overflow_253_fu_24750_p2;
wire   [0:0] xor_ln302_184_fu_24774_p2;
wire   [0:0] underflow_253_fu_24762_p2;
wire   [0:0] or_ln302_91_fu_24780_p2;
wire   [31:0] select_ln302_183_fu_24786_p3;
wire   [31:0] select_ln350_91_fu_24794_p3;
wire  signed [31:0] lhs_74_fu_24006_p3;
wire  signed [31:0] rhs_92_fu_20679_p3;
wire  signed [32:0] sext_ln813_168_fu_24814_p1;
wire  signed [32:0] sext_ln813_167_fu_24810_p1;
wire   [32:0] ret_V_92_fu_24818_p2;
wire   [31:0] p_Val2_669_fu_24832_p2;
wire   [0:0] p_Result_669_fu_24824_p3;
wire   [0:0] p_Result_670_fu_24838_p3;
wire   [0:0] xor_ln895_416_fu_24846_p2;
wire   [0:0] xor_ln896_416_fu_24858_p2;
wire   [0:0] xor_ln302_185_fu_24870_p2;
wire   [0:0] overflow_254_fu_24852_p2;
wire   [0:0] xor_ln302_186_fu_24876_p2;
wire   [0:0] underflow_254_fu_24864_p2;
wire   [0:0] or_ln302_92_fu_24882_p2;
wire   [31:0] select_ln302_185_fu_24888_p3;
wire   [31:0] select_ln350_92_fu_24896_p3;
wire  signed [31:0] lhs_75_fu_24104_p3;
wire  signed [31:0] rhs_93_fu_20828_p3;
wire  signed [32:0] sext_ln813_170_fu_24916_p1;
wire  signed [32:0] sext_ln813_169_fu_24912_p1;
wire   [32:0] ret_V_93_fu_24920_p2;
wire   [31:0] p_Val2_671_fu_24934_p2;
wire   [0:0] p_Result_671_fu_24926_p3;
wire   [0:0] p_Result_672_fu_24940_p3;
wire   [0:0] xor_ln895_417_fu_24948_p2;
wire   [0:0] xor_ln896_417_fu_24960_p2;
wire   [0:0] xor_ln302_187_fu_24972_p2;
wire   [0:0] overflow_255_fu_24954_p2;
wire   [0:0] xor_ln302_188_fu_24978_p2;
wire   [0:0] underflow_255_fu_24966_p2;
wire   [0:0] or_ln302_93_fu_24984_p2;
wire   [31:0] select_ln302_187_fu_24990_p3;
wire   [31:0] select_ln350_93_fu_24998_p3;
wire  signed [31:0] lhs_76_fu_24202_p3;
wire  signed [31:0] rhs_94_fu_20846_p3;
wire  signed [32:0] sext_ln813_172_fu_25018_p1;
wire  signed [32:0] sext_ln813_171_fu_25014_p1;
wire   [32:0] ret_V_94_fu_25022_p2;
wire   [31:0] p_Val2_673_fu_25036_p2;
wire   [0:0] p_Result_673_fu_25028_p3;
wire   [0:0] p_Result_674_fu_25042_p3;
wire   [0:0] xor_ln895_418_fu_25050_p2;
wire   [0:0] xor_ln896_418_fu_25062_p2;
wire   [0:0] xor_ln302_189_fu_25074_p2;
wire   [0:0] overflow_256_fu_25056_p2;
wire   [0:0] xor_ln302_190_fu_25080_p2;
wire   [0:0] underflow_256_fu_25068_p2;
wire   [0:0] or_ln302_94_fu_25086_p2;
wire   [31:0] select_ln302_189_fu_25092_p3;
wire   [31:0] select_ln350_94_fu_25100_p3;
wire  signed [31:0] lhs_77_fu_24300_p3;
wire  signed [31:0] rhs_95_fu_20994_p3;
wire  signed [32:0] sext_ln813_174_fu_25120_p1;
wire  signed [32:0] sext_ln813_173_fu_25116_p1;
wire   [32:0] ret_V_95_fu_25124_p2;
wire   [31:0] p_Val2_675_fu_25138_p2;
wire   [0:0] p_Result_675_fu_25130_p3;
wire   [0:0] p_Result_676_fu_25144_p3;
wire   [0:0] xor_ln895_419_fu_25152_p2;
wire   [0:0] xor_ln896_419_fu_25164_p2;
wire   [0:0] xor_ln302_191_fu_25176_p2;
wire   [0:0] overflow_257_fu_25158_p2;
wire   [0:0] xor_ln302_192_fu_25182_p2;
wire   [0:0] underflow_257_fu_25170_p2;
wire   [0:0] or_ln302_95_fu_25188_p2;
wire   [31:0] select_ln302_191_fu_25194_p3;
wire   [31:0] select_ln350_95_fu_25202_p3;
wire  signed [31:0] lhs_78_fu_24398_p3;
wire  signed [31:0] rhs_96_fu_21143_p3;
wire  signed [32:0] sext_ln813_176_fu_25222_p1;
wire  signed [32:0] sext_ln813_175_fu_25218_p1;
wire   [32:0] ret_V_96_fu_25226_p2;
wire   [31:0] p_Val2_677_fu_25240_p2;
wire   [0:0] p_Result_677_fu_25232_p3;
wire   [0:0] p_Result_678_fu_25246_p3;
wire   [0:0] xor_ln895_420_fu_25254_p2;
wire   [0:0] xor_ln896_420_fu_25266_p2;
wire   [0:0] xor_ln302_193_fu_25278_p2;
wire   [0:0] overflow_258_fu_25260_p2;
wire   [0:0] xor_ln302_194_fu_25284_p2;
wire   [0:0] underflow_258_fu_25272_p2;
wire   [0:0] or_ln302_96_fu_25290_p2;
wire   [31:0] select_ln302_193_fu_25296_p3;
wire   [31:0] select_ln350_96_fu_25304_p3;
wire  signed [31:0] lhs_79_fu_24496_p3;
wire  signed [31:0] rhs_97_fu_21292_p3;
wire  signed [32:0] sext_ln813_178_fu_25324_p1;
wire  signed [32:0] sext_ln813_177_fu_25320_p1;
wire   [32:0] ret_V_97_fu_25328_p2;
wire   [31:0] p_Val2_679_fu_25342_p2;
wire   [0:0] p_Result_679_fu_25334_p3;
wire   [0:0] p_Result_680_fu_25348_p3;
wire   [0:0] xor_ln895_421_fu_25356_p2;
wire   [0:0] xor_ln896_421_fu_25368_p2;
wire   [0:0] xor_ln302_195_fu_25380_p2;
wire   [0:0] overflow_259_fu_25362_p2;
wire   [0:0] xor_ln302_196_fu_25386_p2;
wire   [0:0] underflow_259_fu_25374_p2;
wire   [0:0] or_ln302_97_fu_25392_p2;
wire   [31:0] select_ln302_195_fu_25398_p3;
wire   [31:0] select_ln350_97_fu_25406_p3;
wire   [31:0] select_ln346_181_fu_25425_p3;
wire  signed [31:0] sext_ln856_95_fu_25422_p1;
wire   [31:0] select_ln346_182_fu_25442_p3;
wire  signed [31:0] sext_ln856_96_fu_25439_p1;
wire   [31:0] select_ln346_184_fu_25459_p3;
wire  signed [31:0] sext_ln856_97_fu_25456_p1;
wire   [31:0] select_ln346_185_fu_25476_p3;
wire  signed [31:0] sext_ln856_98_fu_25473_p1;
wire   [31:0] select_ln346_186_fu_25493_p3;
wire  signed [31:0] sext_ln856_99_fu_25490_p1;
wire   [31:0] select_ln346_187_fu_25510_p3;
wire  signed [31:0] sext_ln856_100_fu_25507_p1;
wire   [31:0] select_ln346_188_fu_25527_p3;
wire  signed [31:0] sext_ln856_101_fu_25524_p1;
wire   [0:0] xor_ln896_296_fu_25544_p2;
wire   [0:0] xor_ln888_212_fu_25554_p2;
wire   [0:0] or_ln888_107_fu_25559_p2;
wire   [0:0] tmp_804_fu_25569_p3;
wire   [0:0] xor_ln890_105_fu_25577_p2;
wire   [0:0] or_ln890_107_fu_25583_p2;
wire   [0:0] carry_213_fu_25549_p2;
wire   [0:0] deleted_zeros_104_fu_25564_p2;
wire   [0:0] xor_ln895_296_fu_25599_p2;
wire   [0:0] or_ln895_107_fu_25605_p2;
wire   [0:0] xor_ln895_297_fu_25610_p2;
wire   [0:0] deleted_ones_188_fu_25589_p2;
wire   [0:0] xor_ln896_297_fu_25621_p2;
wire   [0:0] and_ln891_107_fu_25594_p2;
wire   [0:0] or_ln896_107_fu_25627_p2;
wire   [0:0] xor_ln896_512_fu_25633_p2;
wire   [0:0] overflow_188_fu_25615_p2;
wire   [0:0] underflow_188_fu_25639_p2;
wire   [0:0] or_ln346_107_fu_25652_p2;
wire   [31:0] select_ln346_189_fu_25644_p3;
wire  signed [31:0] sext_ln856_102_fu_25541_p1;
wire   [0:0] xor_ln896_298_fu_25669_p2;
wire   [0:0] xor_ln888_214_fu_25679_p2;
wire   [0:0] or_ln888_108_fu_25684_p2;
wire   [0:0] tmp_810_fu_25694_p3;
wire   [0:0] xor_ln890_106_fu_25702_p2;
wire   [0:0] or_ln890_108_fu_25708_p2;
wire   [0:0] carry_215_fu_25674_p2;
wire   [0:0] deleted_zeros_105_fu_25689_p2;
wire   [0:0] xor_ln895_298_fu_25724_p2;
wire   [0:0] or_ln895_108_fu_25730_p2;
wire   [0:0] xor_ln895_299_fu_25735_p2;
wire   [0:0] deleted_ones_189_fu_25714_p2;
wire   [0:0] xor_ln896_299_fu_25746_p2;
wire   [0:0] and_ln891_108_fu_25719_p2;
wire   [0:0] or_ln896_108_fu_25752_p2;
wire   [0:0] xor_ln896_513_fu_25758_p2;
wire   [0:0] overflow_189_fu_25740_p2;
wire   [0:0] underflow_189_fu_25764_p2;
wire   [0:0] or_ln346_108_fu_25777_p2;
wire   [31:0] select_ln346_190_fu_25769_p3;
wire  signed [31:0] sext_ln856_103_fu_25666_p1;
wire   [0:0] xor_ln896_300_fu_25794_p2;
wire   [0:0] xor_ln888_216_fu_25804_p2;
wire   [0:0] or_ln888_109_fu_25809_p2;
wire   [0:0] tmp_816_fu_25819_p3;
wire   [0:0] xor_ln890_107_fu_25827_p2;
wire   [0:0] or_ln890_109_fu_25833_p2;
wire   [0:0] carry_217_fu_25799_p2;
wire   [0:0] deleted_zeros_106_fu_25814_p2;
wire   [0:0] xor_ln895_300_fu_25849_p2;
wire   [0:0] or_ln895_109_fu_25855_p2;
wire   [0:0] xor_ln895_301_fu_25860_p2;
wire   [0:0] deleted_ones_190_fu_25839_p2;
wire   [0:0] xor_ln896_301_fu_25871_p2;
wire   [0:0] and_ln891_109_fu_25844_p2;
wire   [0:0] or_ln896_109_fu_25877_p2;
wire   [0:0] xor_ln896_514_fu_25883_p2;
wire   [0:0] overflow_190_fu_25865_p2;
wire   [0:0] underflow_190_fu_25889_p2;
wire   [0:0] or_ln346_109_fu_25902_p2;
wire   [31:0] select_ln346_191_fu_25894_p3;
wire  signed [31:0] sext_ln856_104_fu_25791_p1;
wire   [0:0] xor_ln896_302_fu_25919_p2;
wire   [0:0] xor_ln888_218_fu_25929_p2;
wire   [0:0] or_ln888_110_fu_25934_p2;
wire   [0:0] tmp_822_fu_25944_p3;
wire   [0:0] xor_ln890_108_fu_25952_p2;
wire   [0:0] or_ln890_110_fu_25958_p2;
wire   [0:0] carry_219_fu_25924_p2;
wire   [0:0] deleted_zeros_107_fu_25939_p2;
wire   [0:0] xor_ln895_302_fu_25974_p2;
wire   [0:0] or_ln895_110_fu_25980_p2;
wire   [0:0] xor_ln895_303_fu_25985_p2;
wire   [0:0] deleted_ones_191_fu_25964_p2;
wire   [0:0] xor_ln896_303_fu_25996_p2;
wire   [0:0] and_ln891_110_fu_25969_p2;
wire   [0:0] or_ln896_110_fu_26002_p2;
wire   [0:0] xor_ln896_515_fu_26008_p2;
wire   [0:0] overflow_191_fu_25990_p2;
wire   [0:0] underflow_191_fu_26014_p2;
wire   [0:0] or_ln346_110_fu_26027_p2;
wire   [31:0] select_ln346_192_fu_26019_p3;
wire  signed [31:0] sext_ln856_105_fu_25916_p1;
wire   [0:0] xor_ln896_304_fu_26044_p2;
wire   [0:0] xor_ln888_220_fu_26054_p2;
wire   [0:0] or_ln888_111_fu_26059_p2;
wire   [0:0] tmp_828_fu_26069_p3;
wire   [0:0] xor_ln890_109_fu_26077_p2;
wire   [0:0] or_ln890_111_fu_26083_p2;
wire   [0:0] carry_221_fu_26049_p2;
wire   [0:0] deleted_zeros_108_fu_26064_p2;
wire   [0:0] xor_ln895_304_fu_26099_p2;
wire   [0:0] or_ln895_111_fu_26105_p2;
wire   [0:0] xor_ln895_305_fu_26110_p2;
wire   [0:0] deleted_ones_192_fu_26089_p2;
wire   [0:0] xor_ln896_305_fu_26121_p2;
wire   [0:0] and_ln891_111_fu_26094_p2;
wire   [0:0] or_ln896_111_fu_26127_p2;
wire   [0:0] xor_ln896_516_fu_26133_p2;
wire   [0:0] overflow_192_fu_26115_p2;
wire   [0:0] underflow_192_fu_26139_p2;
wire   [0:0] or_ln346_111_fu_26152_p2;
wire   [31:0] select_ln346_193_fu_26144_p3;
wire  signed [31:0] sext_ln856_106_fu_26041_p1;
wire   [0:0] xor_ln896_306_fu_26169_p2;
wire   [0:0] xor_ln888_222_fu_26179_p2;
wire   [0:0] or_ln888_112_fu_26184_p2;
wire   [0:0] tmp_834_fu_26194_p3;
wire   [0:0] xor_ln890_110_fu_26202_p2;
wire   [0:0] or_ln890_112_fu_26208_p2;
wire   [0:0] carry_223_fu_26174_p2;
wire   [0:0] deleted_zeros_109_fu_26189_p2;
wire   [0:0] xor_ln895_306_fu_26224_p2;
wire   [0:0] or_ln895_112_fu_26230_p2;
wire   [0:0] xor_ln895_307_fu_26235_p2;
wire   [0:0] deleted_ones_193_fu_26214_p2;
wire   [0:0] xor_ln896_307_fu_26246_p2;
wire   [0:0] and_ln891_112_fu_26219_p2;
wire   [0:0] or_ln896_112_fu_26252_p2;
wire   [0:0] xor_ln896_517_fu_26258_p2;
wire   [0:0] overflow_193_fu_26240_p2;
wire   [0:0] underflow_193_fu_26264_p2;
wire   [0:0] or_ln346_112_fu_26277_p2;
wire   [31:0] select_ln346_194_fu_26269_p3;
wire  signed [31:0] sext_ln856_107_fu_26166_p1;
wire   [31:0] select_ln346_195_fu_26294_p3;
wire  signed [31:0] sext_ln856_108_fu_26291_p1;
wire   [0:0] xor_ln896_310_fu_26311_p2;
wire   [0:0] xor_ln888_226_fu_26321_p2;
wire   [0:0] or_ln888_114_fu_26326_p2;
wire   [0:0] tmp_846_fu_26336_p3;
wire   [0:0] xor_ln890_112_fu_26344_p2;
wire   [0:0] or_ln890_114_fu_26350_p2;
wire   [0:0] carry_227_fu_26316_p2;
wire   [0:0] deleted_zeros_111_fu_26331_p2;
wire   [0:0] xor_ln895_310_fu_26366_p2;
wire   [0:0] or_ln895_114_fu_26372_p2;
wire   [0:0] xor_ln895_311_fu_26377_p2;
wire   [0:0] deleted_ones_195_fu_26356_p2;
wire   [0:0] xor_ln896_311_fu_26388_p2;
wire   [0:0] and_ln891_114_fu_26361_p2;
wire   [0:0] or_ln896_114_fu_26394_p2;
wire   [0:0] xor_ln896_519_fu_26400_p2;
wire   [0:0] overflow_195_fu_26382_p2;
wire   [0:0] underflow_195_fu_26406_p2;
wire   [0:0] or_ln346_114_fu_26419_p2;
wire   [31:0] select_ln346_196_fu_26411_p3;
wire  signed [31:0] sext_ln856_109_fu_26308_p1;
wire   [0:0] xor_ln896_312_fu_26436_p2;
wire   [0:0] xor_ln888_228_fu_26446_p2;
wire   [0:0] or_ln888_115_fu_26451_p2;
wire   [0:0] tmp_852_fu_26461_p3;
wire   [0:0] xor_ln890_113_fu_26469_p2;
wire   [0:0] or_ln890_115_fu_26475_p2;
wire   [0:0] carry_229_fu_26441_p2;
wire   [0:0] deleted_zeros_112_fu_26456_p2;
wire   [0:0] xor_ln895_312_fu_26491_p2;
wire   [0:0] or_ln895_115_fu_26497_p2;
wire   [0:0] xor_ln895_313_fu_26502_p2;
wire   [0:0] deleted_ones_196_fu_26481_p2;
wire   [0:0] xor_ln896_313_fu_26513_p2;
wire   [0:0] and_ln891_115_fu_26486_p2;
wire   [0:0] or_ln896_115_fu_26519_p2;
wire   [0:0] xor_ln896_520_fu_26525_p2;
wire   [0:0] overflow_196_fu_26507_p2;
wire   [0:0] underflow_196_fu_26531_p2;
wire   [0:0] or_ln346_115_fu_26544_p2;
wire   [31:0] select_ln346_197_fu_26536_p3;
wire  signed [31:0] sext_ln856_110_fu_26433_p1;
wire   [31:0] zext_ln377_116_fu_26561_p1;
wire  signed [31:0] sext_ln818_1_fu_26558_p1;
wire   [31:0] p_Val2_511_fu_26564_p2;
wire   [0:0] p_Result_512_fu_26570_p3;
wire   [0:0] xor_ln896_314_fu_26578_p2;
wire   [0:0] xor_ln888_230_fu_26589_p2;
wire   [0:0] or_ln888_116_fu_26594_p2;
wire   [0:0] tmp_858_fu_26605_p3;
wire   [0:0] xor_ln890_114_fu_26613_p2;
wire   [0:0] or_ln890_116_fu_26619_p2;
wire   [0:0] carry_231_fu_26584_p2;
wire   [0:0] deleted_zeros_113_fu_26600_p2;
wire   [0:0] xor_ln895_314_fu_26635_p2;
wire   [0:0] or_ln895_116_fu_26641_p2;
wire   [0:0] xor_ln895_315_fu_26647_p2;
wire   [0:0] deleted_ones_197_fu_26625_p2;
wire   [0:0] xor_ln896_315_fu_26658_p2;
wire   [0:0] and_ln891_116_fu_26630_p2;
wire   [0:0] or_ln896_116_fu_26664_p2;
wire   [0:0] xor_ln896_521_fu_26670_p2;
wire   [0:0] overflow_197_fu_26652_p2;
wire   [0:0] underflow_197_fu_26676_p2;
wire   [0:0] or_ln346_116_fu_26689_p2;
wire   [31:0] select_ln346_198_fu_26681_p3;
wire   [18:0] zext_ln377_117_fu_26706_p1;
wire  signed [18:0] sext_ln823_111_fu_26703_p1;
wire  signed [18:0] p_Val2_514_fu_26709_p2;
wire   [0:0] p_Result_515_fu_26719_p3;
wire   [0:0] xor_ln896_316_fu_26727_p2;
wire   [0:0] xor_ln888_232_fu_26738_p2;
wire   [0:0] or_ln888_117_fu_26743_p2;
wire   [0:0] tmp_864_fu_26754_p3;
wire   [0:0] xor_ln890_115_fu_26762_p2;
wire   [0:0] or_ln890_117_fu_26768_p2;
wire   [0:0] carry_233_fu_26733_p2;
wire   [0:0] deleted_zeros_114_fu_26749_p2;
wire   [0:0] xor_ln895_316_fu_26784_p2;
wire   [0:0] or_ln895_117_fu_26790_p2;
wire   [0:0] xor_ln895_317_fu_26796_p2;
wire   [0:0] deleted_ones_198_fu_26774_p2;
wire   [0:0] xor_ln896_317_fu_26807_p2;
wire   [0:0] and_ln891_117_fu_26779_p2;
wire   [0:0] or_ln896_117_fu_26813_p2;
wire   [0:0] xor_ln896_522_fu_26819_p2;
wire   [0:0] overflow_198_fu_26801_p2;
wire   [0:0] underflow_198_fu_26825_p2;
wire   [0:0] or_ln346_117_fu_26838_p2;
wire   [31:0] select_ln346_199_fu_26830_p3;
wire  signed [31:0] sext_ln856_111_fu_26715_p1;
wire   [21:0] zext_ln377_118_fu_26855_p1;
wire  signed [21:0] sext_ln823_112_fu_26852_p1;
wire  signed [21:0] p_Val2_517_fu_26858_p2;
wire   [0:0] p_Result_518_fu_26868_p3;
wire   [0:0] xor_ln896_318_fu_26876_p2;
wire   [0:0] xor_ln888_234_fu_26887_p2;
wire   [0:0] or_ln888_118_fu_26892_p2;
wire   [0:0] tmp_870_fu_26903_p3;
wire   [0:0] xor_ln890_116_fu_26911_p2;
wire   [0:0] or_ln890_118_fu_26917_p2;
wire   [0:0] carry_235_fu_26882_p2;
wire   [0:0] deleted_zeros_115_fu_26898_p2;
wire   [0:0] xor_ln895_318_fu_26933_p2;
wire   [0:0] or_ln895_118_fu_26939_p2;
wire   [0:0] xor_ln895_319_fu_26945_p2;
wire   [0:0] deleted_ones_199_fu_26923_p2;
wire   [0:0] xor_ln896_319_fu_26956_p2;
wire   [0:0] and_ln891_118_fu_26928_p2;
wire   [0:0] or_ln896_118_fu_26962_p2;
wire   [0:0] xor_ln896_523_fu_26968_p2;
wire   [0:0] overflow_199_fu_26950_p2;
wire   [0:0] underflow_199_fu_26974_p2;
wire   [0:0] or_ln346_118_fu_26987_p2;
wire   [31:0] select_ln346_200_fu_26979_p3;
wire  signed [31:0] sext_ln856_112_fu_26864_p1;
wire   [21:0] zext_ln377_119_fu_27004_p1;
wire  signed [21:0] sext_ln823_113_fu_27001_p1;
wire  signed [21:0] p_Val2_520_fu_27007_p2;
wire   [0:0] p_Result_521_fu_27017_p3;
wire   [0:0] xor_ln896_320_fu_27025_p2;
wire   [0:0] xor_ln888_236_fu_27036_p2;
wire   [0:0] or_ln888_119_fu_27041_p2;
wire   [0:0] tmp_876_fu_27052_p3;
wire   [0:0] xor_ln890_117_fu_27060_p2;
wire   [0:0] or_ln890_119_fu_27066_p2;
wire   [0:0] carry_237_fu_27031_p2;
wire   [0:0] deleted_zeros_116_fu_27047_p2;
wire   [0:0] xor_ln895_320_fu_27082_p2;
wire   [0:0] or_ln895_119_fu_27088_p2;
wire   [0:0] xor_ln895_321_fu_27094_p2;
wire   [0:0] deleted_ones_200_fu_27072_p2;
wire   [0:0] xor_ln896_321_fu_27105_p2;
wire   [0:0] and_ln891_119_fu_27077_p2;
wire   [0:0] or_ln896_119_fu_27111_p2;
wire   [0:0] xor_ln896_524_fu_27117_p2;
wire   [0:0] overflow_200_fu_27099_p2;
wire   [0:0] underflow_200_fu_27123_p2;
wire   [0:0] or_ln346_119_fu_27136_p2;
wire   [31:0] select_ln346_201_fu_27128_p3;
wire  signed [31:0] sext_ln856_113_fu_27013_p1;
wire   [23:0] zext_ln377_120_fu_27153_p1;
wire  signed [23:0] sext_ln823_114_fu_27150_p1;
wire  signed [23:0] p_Val2_523_fu_27156_p2;
wire   [0:0] p_Result_524_fu_27166_p3;
wire   [0:0] xor_ln896_322_fu_27174_p2;
wire   [0:0] xor_ln888_238_fu_27185_p2;
wire   [0:0] or_ln888_120_fu_27190_p2;
wire   [0:0] tmp_882_fu_27201_p3;
wire   [0:0] xor_ln890_118_fu_27209_p2;
wire   [0:0] or_ln890_120_fu_27215_p2;
wire   [0:0] carry_239_fu_27180_p2;
wire   [0:0] deleted_zeros_117_fu_27196_p2;
wire   [0:0] xor_ln895_322_fu_27231_p2;
wire   [0:0] or_ln895_120_fu_27237_p2;
wire   [0:0] xor_ln895_323_fu_27243_p2;
wire   [0:0] deleted_ones_201_fu_27221_p2;
wire   [0:0] xor_ln896_323_fu_27254_p2;
wire   [0:0] and_ln891_120_fu_27226_p2;
wire   [0:0] or_ln896_120_fu_27260_p2;
wire   [0:0] xor_ln896_525_fu_27266_p2;
wire   [0:0] overflow_201_fu_27248_p2;
wire   [0:0] underflow_201_fu_27272_p2;
wire   [0:0] or_ln346_120_fu_27285_p2;
wire   [31:0] select_ln346_202_fu_27277_p3;
wire  signed [31:0] sext_ln856_114_fu_27162_p1;
wire   [19:0] zext_ln377_121_fu_27302_p1;
wire  signed [19:0] sext_ln823_115_fu_27299_p1;
wire  signed [19:0] p_Val2_526_fu_27305_p2;
wire   [0:0] p_Result_527_fu_27315_p3;
wire   [0:0] xor_ln896_324_fu_27323_p2;
wire   [0:0] xor_ln888_240_fu_27334_p2;
wire   [0:0] or_ln888_121_fu_27339_p2;
wire   [0:0] tmp_888_fu_27350_p3;
wire   [0:0] xor_ln890_119_fu_27358_p2;
wire   [0:0] or_ln890_121_fu_27364_p2;
wire   [0:0] carry_241_fu_27329_p2;
wire   [0:0] deleted_zeros_118_fu_27345_p2;
wire   [0:0] xor_ln895_324_fu_27380_p2;
wire   [0:0] or_ln895_121_fu_27386_p2;
wire   [0:0] xor_ln895_325_fu_27392_p2;
wire   [0:0] deleted_ones_202_fu_27370_p2;
wire   [0:0] xor_ln896_325_fu_27403_p2;
wire   [0:0] and_ln891_121_fu_27375_p2;
wire   [0:0] or_ln896_121_fu_27409_p2;
wire   [0:0] xor_ln896_526_fu_27415_p2;
wire   [0:0] overflow_202_fu_27397_p2;
wire   [0:0] underflow_202_fu_27421_p2;
wire   [0:0] or_ln346_121_fu_27434_p2;
wire   [31:0] select_ln346_203_fu_27426_p3;
wire  signed [31:0] sext_ln856_115_fu_27311_p1;
wire   [21:0] zext_ln377_122_fu_27451_p1;
wire  signed [21:0] sext_ln823_116_fu_27448_p1;
wire  signed [21:0] p_Val2_529_fu_27454_p2;
wire   [0:0] p_Result_530_fu_27464_p3;
wire   [0:0] xor_ln896_326_fu_27472_p2;
wire   [0:0] xor_ln888_242_fu_27483_p2;
wire   [0:0] or_ln888_122_fu_27488_p2;
wire   [0:0] tmp_894_fu_27499_p3;
wire   [0:0] xor_ln890_120_fu_27507_p2;
wire   [0:0] or_ln890_122_fu_27513_p2;
wire   [0:0] carry_243_fu_27478_p2;
wire   [0:0] deleted_zeros_119_fu_27494_p2;
wire   [0:0] xor_ln895_326_fu_27529_p2;
wire   [0:0] or_ln895_122_fu_27535_p2;
wire   [0:0] xor_ln895_327_fu_27541_p2;
wire   [0:0] deleted_ones_203_fu_27519_p2;
wire   [0:0] xor_ln896_327_fu_27552_p2;
wire   [0:0] and_ln891_122_fu_27524_p2;
wire   [0:0] or_ln896_122_fu_27558_p2;
wire   [0:0] xor_ln896_527_fu_27564_p2;
wire   [0:0] overflow_203_fu_27546_p2;
wire   [0:0] underflow_203_fu_27570_p2;
wire   [0:0] or_ln346_122_fu_27583_p2;
wire   [31:0] select_ln346_204_fu_27575_p3;
wire  signed [31:0] sext_ln856_116_fu_27460_p1;
wire   [20:0] zext_ln377_123_fu_27600_p1;
wire  signed [20:0] sext_ln823_117_fu_27597_p1;
wire  signed [20:0] p_Val2_532_fu_27603_p2;
wire   [0:0] p_Result_533_fu_27613_p3;
wire   [0:0] xor_ln896_328_fu_27621_p2;
wire   [0:0] xor_ln888_244_fu_27632_p2;
wire   [0:0] or_ln888_123_fu_27637_p2;
wire   [0:0] tmp_900_fu_27648_p3;
wire   [0:0] xor_ln890_121_fu_27656_p2;
wire   [0:0] or_ln890_123_fu_27662_p2;
wire   [0:0] carry_245_fu_27627_p2;
wire   [0:0] deleted_zeros_120_fu_27643_p2;
wire   [0:0] xor_ln895_328_fu_27678_p2;
wire   [0:0] or_ln895_123_fu_27684_p2;
wire   [0:0] xor_ln895_329_fu_27690_p2;
wire   [0:0] deleted_ones_204_fu_27668_p2;
wire   [0:0] xor_ln896_329_fu_27701_p2;
wire   [0:0] and_ln891_123_fu_27673_p2;
wire   [0:0] or_ln896_123_fu_27707_p2;
wire   [0:0] xor_ln896_528_fu_27713_p2;
wire   [0:0] overflow_204_fu_27695_p2;
wire   [0:0] underflow_204_fu_27719_p2;
wire   [0:0] or_ln346_123_fu_27732_p2;
wire   [31:0] select_ln346_205_fu_27724_p3;
wire  signed [31:0] sext_ln856_117_fu_27609_p1;
wire   [20:0] zext_ln377_124_fu_27749_p1;
wire  signed [20:0] sext_ln823_118_fu_27746_p1;
wire  signed [20:0] p_Val2_535_fu_27752_p2;
wire   [0:0] p_Result_536_fu_27762_p3;
wire   [0:0] xor_ln896_330_fu_27770_p2;
wire   [0:0] xor_ln888_246_fu_27781_p2;
wire   [0:0] or_ln888_124_fu_27786_p2;
wire   [0:0] tmp_906_fu_27797_p3;
wire   [0:0] xor_ln890_122_fu_27805_p2;
wire   [0:0] or_ln890_124_fu_27811_p2;
wire   [0:0] carry_247_fu_27776_p2;
wire   [0:0] deleted_zeros_121_fu_27792_p2;
wire   [0:0] xor_ln895_330_fu_27827_p2;
wire   [0:0] or_ln895_124_fu_27833_p2;
wire   [0:0] xor_ln895_331_fu_27839_p2;
wire   [0:0] deleted_ones_205_fu_27817_p2;
wire   [0:0] xor_ln896_331_fu_27850_p2;
wire   [0:0] and_ln891_124_fu_27822_p2;
wire   [0:0] or_ln896_124_fu_27856_p2;
wire   [0:0] xor_ln896_529_fu_27862_p2;
wire   [0:0] overflow_205_fu_27844_p2;
wire   [0:0] underflow_205_fu_27868_p2;
wire   [0:0] or_ln346_124_fu_27881_p2;
wire   [31:0] select_ln346_206_fu_27873_p3;
wire  signed [31:0] sext_ln856_118_fu_27758_p1;
wire   [39:0] shl_ln1273_14_fu_27918_p3;
wire   [32:0] shl_ln1273_15_fu_27929_p3;
wire  signed [40:0] sext_ln1273_17_fu_27936_p1;
wire  signed [40:0] sext_ln1273_16_fu_27925_p1;
wire   [40:0] r_V_122_fu_27940_p2;
wire   [16:0] p_Val2_537_fu_27954_p4;
wire   [17:0] zext_ln377_125_fu_27976_p1;
wire  signed [17:0] sext_ln823_119_fu_27964_p1;
wire   [0:0] p_Result_539_fu_27985_p3;
wire   [0:0] p_Result_538_fu_27968_p3;
wire   [0:0] xor_ln896_332_fu_27993_p2;
wire   [0:0] xor_ln888_248_fu_28013_p2;
wire   [0:0] Range2_all_ones_123_fu_28005_p3;
wire   [0:0] or_ln888_125_fu_28019_p2;
wire   [0:0] tmp_912_fu_28031_p3;
wire   [0:0] xor_ln890_123_fu_28039_p2;
wire   [0:0] or_ln890_125_fu_28045_p2;
wire   [0:0] carry_249_fu_27999_p2;
wire   [0:0] deleted_zeros_122_fu_28025_p2;
wire   [0:0] xor_ln895_332_fu_28063_p2;
wire   [0:0] p_Result_537_fu_27946_p3;
wire   [0:0] or_ln895_125_fu_28069_p2;
wire   [0:0] xor_ln895_333_fu_28075_p2;
wire   [0:0] deleted_ones_206_fu_28051_p2;
wire   [0:0] xor_ln896_333_fu_28087_p2;
wire   [0:0] and_ln891_125_fu_28057_p2;
wire   [0:0] or_ln896_125_fu_28093_p2;
wire   [0:0] xor_ln896_530_fu_28099_p2;
wire   [0:0] underflow_206_fu_28105_p2;
wire   [18:0] p_Val2_540_fu_28125_p4;
wire   [0:0] tmp_915_fu_28147_p3;
wire   [19:0] zext_ln377_126_fu_28155_p1;
wire  signed [19:0] sext_ln823_120_fu_28135_p1;
wire   [19:0] p_Val2_543_fu_28189_p4;
wire   [0:0] tmp_921_fu_28211_p3;
wire   [20:0] zext_ln377_127_fu_28219_p1;
wire  signed [20:0] sext_ln823_121_fu_28199_p1;
wire   [18:0] p_Val2_546_fu_28253_p4;
wire   [0:0] tmp_927_fu_28275_p3;
wire   [19:0] zext_ln377_128_fu_28283_p1;
wire  signed [19:0] sext_ln823_122_fu_28263_p1;
wire   [19:0] p_Val2_549_fu_28317_p4;
wire   [0:0] tmp_933_fu_28339_p3;
wire   [20:0] zext_ln377_129_fu_28347_p1;
wire  signed [20:0] sext_ln823_123_fu_28327_p1;
wire   [18:0] p_Val2_552_fu_28381_p4;
wire   [0:0] tmp_939_fu_28403_p3;
wire   [19:0] zext_ln377_130_fu_28411_p1;
wire  signed [19:0] sext_ln823_124_fu_28391_p1;
wire   [20:0] p_Val2_555_fu_28445_p4;
wire   [0:0] tmp_945_fu_28467_p3;
wire   [21:0] zext_ln377_131_fu_28475_p1;
wire  signed [21:0] sext_ln823_125_fu_28455_p1;
wire   [15:0] p_Val2_558_fu_28509_p4;
wire   [0:0] tmp_951_fu_28531_p3;
wire   [16:0] zext_ln377_132_fu_28539_p1;
wire  signed [16:0] sext_ln823_126_fu_28519_p1;
wire   [17:0] p_Val2_561_fu_28573_p4;
wire   [0:0] tmp_957_fu_28595_p3;
wire   [18:0] zext_ln377_133_fu_28603_p1;
wire  signed [18:0] sext_ln823_127_fu_28583_p1;
wire   [39:0] shl_ln1273_16_fu_28985_p3;
wire   [36:0] shl_ln1273_17_fu_28996_p3;
wire  signed [40:0] sext_ln1273_19_fu_29003_p1;
wire  signed [40:0] sext_ln1273_18_fu_28992_p1;
wire   [40:0] r_V_139_fu_29007_p2;
wire   [16:0] p_Val2_588_fu_29021_p4;
wire   [17:0] zext_ln377_142_fu_29043_p1;
wire  signed [17:0] sext_ln823_136_fu_29031_p1;
wire   [0:0] p_Result_590_fu_29052_p3;
wire   [0:0] p_Result_589_fu_29035_p3;
wire   [0:0] xor_ln896_366_fu_29060_p2;
wire   [0:0] xor_ln888_282_fu_29080_p2;
wire   [0:0] Range2_all_ones_140_fu_29072_p3;
wire   [0:0] or_ln888_142_fu_29086_p2;
wire   [0:0] tmp_1014_fu_29098_p3;
wire   [0:0] xor_ln890_140_fu_29106_p2;
wire   [0:0] or_ln890_142_fu_29112_p2;
wire   [0:0] carry_283_fu_29066_p2;
wire   [0:0] deleted_zeros_139_fu_29092_p2;
wire   [0:0] xor_ln895_366_fu_29130_p2;
wire   [0:0] p_Result_588_fu_29013_p3;
wire   [0:0] or_ln895_142_fu_29136_p2;
wire   [0:0] xor_ln895_367_fu_29142_p2;
wire   [0:0] deleted_ones_223_fu_29118_p2;
wire   [0:0] xor_ln896_367_fu_29154_p2;
wire   [0:0] and_ln891_142_fu_29124_p2;
wire   [0:0] or_ln896_142_fu_29160_p2;
wire   [0:0] xor_ln896_547_fu_29166_p2;
wire   [0:0] underflow_223_fu_29172_p2;
wire  signed [32:0] sext_ln813_180_fu_29187_p1;
wire  signed [32:0] sext_ln813_179_fu_29184_p1;
wire   [32:0] ret_V_98_fu_29190_p2;
wire   [31:0] p_Val2_681_fu_29204_p2;
wire   [0:0] p_Result_681_fu_29196_p3;
wire   [0:0] p_Result_682_fu_29208_p3;
wire   [0:0] xor_ln895_422_fu_29216_p2;
wire   [0:0] xor_ln896_422_fu_29228_p2;
wire   [0:0] xor_ln302_197_fu_29240_p2;
wire   [0:0] overflow_260_fu_29222_p2;
wire   [0:0] xor_ln302_198_fu_29246_p2;
wire   [0:0] underflow_260_fu_29234_p2;
wire   [0:0] or_ln302_98_fu_29252_p2;
wire   [31:0] select_ln302_197_fu_29258_p3;
wire   [31:0] select_ln350_98_fu_29266_p3;
wire  signed [31:0] rhs_99_fu_25432_p3;
wire  signed [32:0] sext_ln813_182_fu_29285_p1;
wire  signed [32:0] sext_ln813_181_fu_29282_p1;
wire   [32:0] ret_V_99_fu_29289_p2;
wire   [31:0] p_Val2_683_fu_29303_p2;
wire   [0:0] p_Result_683_fu_29295_p3;
wire   [0:0] p_Result_684_fu_29308_p3;
wire   [0:0] xor_ln895_423_fu_29316_p2;
wire   [0:0] xor_ln896_423_fu_29328_p2;
wire   [0:0] xor_ln302_199_fu_29340_p2;
wire   [0:0] overflow_261_fu_29322_p2;
wire   [0:0] xor_ln302_200_fu_29346_p2;
wire   [0:0] underflow_261_fu_29334_p2;
wire   [0:0] or_ln302_99_fu_29352_p2;
wire   [31:0] select_ln302_199_fu_29358_p3;
wire   [31:0] select_ln350_99_fu_29366_p3;
wire  signed [31:0] rhs_100_fu_25449_p3;
wire  signed [32:0] sext_ln813_184_fu_29385_p1;
wire  signed [32:0] sext_ln813_183_fu_29382_p1;
wire   [32:0] ret_V_100_fu_29389_p2;
wire   [31:0] p_Val2_685_fu_29403_p2;
wire   [0:0] p_Result_685_fu_29395_p3;
wire   [0:0] p_Result_686_fu_29408_p3;
wire   [0:0] xor_ln895_424_fu_29416_p2;
wire   [0:0] xor_ln896_424_fu_29428_p2;
wire   [0:0] xor_ln302_201_fu_29440_p2;
wire   [0:0] overflow_262_fu_29422_p2;
wire   [0:0] xor_ln302_202_fu_29446_p2;
wire   [0:0] underflow_262_fu_29434_p2;
wire   [0:0] or_ln302_100_fu_29452_p2;
wire   [31:0] select_ln302_201_fu_29458_p3;
wire   [31:0] select_ln350_100_fu_29466_p3;
wire  signed [32:0] sext_ln813_186_fu_29485_p1;
wire  signed [32:0] sext_ln813_185_fu_29482_p1;
wire   [32:0] ret_V_101_fu_29488_p2;
wire   [31:0] p_Val2_687_fu_29502_p2;
wire   [0:0] p_Result_687_fu_29494_p3;
wire   [0:0] p_Result_688_fu_29506_p3;
wire   [0:0] xor_ln895_425_fu_29514_p2;
wire   [0:0] xor_ln896_425_fu_29526_p2;
wire   [0:0] xor_ln302_203_fu_29538_p2;
wire   [0:0] overflow_263_fu_29520_p2;
wire   [0:0] xor_ln302_204_fu_29544_p2;
wire   [0:0] underflow_263_fu_29532_p2;
wire   [0:0] or_ln302_101_fu_29550_p2;
wire   [31:0] select_ln302_203_fu_29556_p3;
wire   [31:0] select_ln350_101_fu_29564_p3;
wire  signed [31:0] rhs_102_fu_25466_p3;
wire  signed [32:0] sext_ln813_188_fu_29583_p1;
wire  signed [32:0] sext_ln813_187_fu_29580_p1;
wire   [32:0] ret_V_102_fu_29587_p2;
wire   [31:0] p_Val2_689_fu_29601_p2;
wire   [0:0] p_Result_689_fu_29593_p3;
wire   [0:0] p_Result_690_fu_29606_p3;
wire   [0:0] xor_ln895_426_fu_29614_p2;
wire   [0:0] xor_ln896_426_fu_29626_p2;
wire   [0:0] xor_ln302_205_fu_29638_p2;
wire   [0:0] overflow_264_fu_29620_p2;
wire   [0:0] xor_ln302_206_fu_29644_p2;
wire   [0:0] underflow_264_fu_29632_p2;
wire   [0:0] or_ln302_102_fu_29650_p2;
wire   [31:0] select_ln302_205_fu_29656_p3;
wire   [31:0] select_ln350_102_fu_29664_p3;
wire  signed [31:0] rhs_103_fu_25483_p3;
wire  signed [32:0] sext_ln813_190_fu_29683_p1;
wire  signed [32:0] sext_ln813_189_fu_29680_p1;
wire   [32:0] ret_V_103_fu_29687_p2;
wire   [31:0] p_Val2_691_fu_29701_p2;
wire   [0:0] p_Result_691_fu_29693_p3;
wire   [0:0] p_Result_692_fu_29706_p3;
wire   [0:0] xor_ln895_427_fu_29714_p2;
wire   [0:0] xor_ln896_427_fu_29726_p2;
wire   [0:0] xor_ln302_207_fu_29738_p2;
wire   [0:0] overflow_265_fu_29720_p2;
wire   [0:0] xor_ln302_208_fu_29744_p2;
wire   [0:0] underflow_265_fu_29732_p2;
wire   [0:0] or_ln302_103_fu_29750_p2;
wire   [31:0] select_ln302_207_fu_29756_p3;
wire   [31:0] select_ln350_103_fu_29764_p3;
wire  signed [31:0] rhs_104_fu_25500_p3;
wire  signed [32:0] sext_ln813_192_fu_29783_p1;
wire  signed [32:0] sext_ln813_191_fu_29780_p1;
wire   [32:0] ret_V_104_fu_29787_p2;
wire   [31:0] p_Val2_693_fu_29801_p2;
wire   [0:0] p_Result_693_fu_29793_p3;
wire   [0:0] p_Result_694_fu_29806_p3;
wire   [0:0] xor_ln895_428_fu_29814_p2;
wire   [0:0] xor_ln896_428_fu_29826_p2;
wire   [0:0] xor_ln302_209_fu_29838_p2;
wire   [0:0] overflow_266_fu_29820_p2;
wire   [0:0] xor_ln302_210_fu_29844_p2;
wire   [0:0] underflow_266_fu_29832_p2;
wire   [0:0] or_ln302_104_fu_29850_p2;
wire   [31:0] select_ln302_209_fu_29856_p3;
wire   [31:0] select_ln350_104_fu_29864_p3;
wire  signed [31:0] rhs_105_fu_25517_p3;
wire  signed [32:0] sext_ln813_194_fu_29883_p1;
wire  signed [32:0] sext_ln813_193_fu_29880_p1;
wire   [32:0] ret_V_105_fu_29887_p2;
wire   [31:0] p_Val2_695_fu_29901_p2;
wire   [0:0] p_Result_695_fu_29893_p3;
wire   [0:0] p_Result_696_fu_29906_p3;
wire   [0:0] xor_ln895_429_fu_29914_p2;
wire   [0:0] xor_ln896_429_fu_29926_p2;
wire   [0:0] xor_ln302_211_fu_29938_p2;
wire   [0:0] overflow_267_fu_29920_p2;
wire   [0:0] xor_ln302_212_fu_29944_p2;
wire   [0:0] underflow_267_fu_29932_p2;
wire   [0:0] or_ln302_105_fu_29950_p2;
wire   [31:0] select_ln302_211_fu_29956_p3;
wire   [31:0] select_ln350_105_fu_29964_p3;
wire  signed [31:0] rhs_106_fu_25534_p3;
wire  signed [32:0] sext_ln813_196_fu_29983_p1;
wire  signed [32:0] sext_ln813_195_fu_29980_p1;
wire   [32:0] ret_V_106_fu_29987_p2;
wire   [31:0] p_Val2_697_fu_30001_p2;
wire   [0:0] p_Result_697_fu_29993_p3;
wire   [0:0] p_Result_698_fu_30006_p3;
wire   [0:0] xor_ln895_430_fu_30014_p2;
wire   [0:0] xor_ln896_430_fu_30026_p2;
wire   [0:0] xor_ln302_213_fu_30038_p2;
wire   [0:0] overflow_268_fu_30020_p2;
wire   [0:0] xor_ln302_214_fu_30044_p2;
wire   [0:0] underflow_268_fu_30032_p2;
wire   [0:0] or_ln302_106_fu_30050_p2;
wire   [31:0] select_ln302_213_fu_30056_p3;
wire   [31:0] select_ln350_106_fu_30064_p3;
wire  signed [31:0] lhs_89_fu_29274_p3;
wire  signed [31:0] rhs_107_fu_25658_p3;
wire  signed [32:0] sext_ln813_198_fu_30084_p1;
wire  signed [32:0] sext_ln813_197_fu_30080_p1;
wire   [32:0] ret_V_107_fu_30088_p2;
wire   [31:0] p_Val2_699_fu_30102_p2;
wire   [0:0] p_Result_699_fu_30094_p3;
wire   [0:0] p_Result_700_fu_30108_p3;
wire   [0:0] xor_ln895_431_fu_30116_p2;
wire   [0:0] xor_ln896_431_fu_30128_p2;
wire   [0:0] xor_ln302_215_fu_30140_p2;
wire   [0:0] overflow_269_fu_30122_p2;
wire   [0:0] xor_ln302_216_fu_30146_p2;
wire   [0:0] underflow_269_fu_30134_p2;
wire   [0:0] or_ln302_107_fu_30152_p2;
wire   [31:0] select_ln302_215_fu_30158_p3;
wire   [31:0] select_ln350_107_fu_30166_p3;
wire  signed [31:0] lhs_90_fu_29374_p3;
wire  signed [31:0] rhs_108_fu_25783_p3;
wire  signed [32:0] sext_ln813_200_fu_30186_p1;
wire  signed [32:0] sext_ln813_199_fu_30182_p1;
wire   [32:0] ret_V_108_fu_30190_p2;
wire   [31:0] p_Val2_701_fu_30204_p2;
wire   [0:0] p_Result_701_fu_30196_p3;
wire   [0:0] p_Result_702_fu_30210_p3;
wire   [0:0] xor_ln895_432_fu_30218_p2;
wire   [0:0] xor_ln896_432_fu_30230_p2;
wire   [0:0] xor_ln302_217_fu_30242_p2;
wire   [0:0] overflow_270_fu_30224_p2;
wire   [0:0] xor_ln302_218_fu_30248_p2;
wire   [0:0] underflow_270_fu_30236_p2;
wire   [0:0] or_ln302_108_fu_30254_p2;
wire   [31:0] select_ln302_217_fu_30260_p3;
wire   [31:0] select_ln350_108_fu_30268_p3;
wire  signed [31:0] lhs_91_fu_29474_p3;
wire  signed [31:0] rhs_109_fu_25908_p3;
wire  signed [32:0] sext_ln813_202_fu_30288_p1;
wire  signed [32:0] sext_ln813_201_fu_30284_p1;
wire   [32:0] ret_V_109_fu_30292_p2;
wire   [31:0] p_Val2_703_fu_30306_p2;
wire   [0:0] p_Result_703_fu_30298_p3;
wire   [0:0] p_Result_704_fu_30312_p3;
wire   [0:0] xor_ln895_433_fu_30320_p2;
wire   [0:0] xor_ln896_433_fu_30332_p2;
wire   [0:0] xor_ln302_219_fu_30344_p2;
wire   [0:0] overflow_271_fu_30326_p2;
wire   [0:0] xor_ln302_220_fu_30350_p2;
wire   [0:0] underflow_271_fu_30338_p2;
wire   [0:0] or_ln302_109_fu_30356_p2;
wire   [31:0] select_ln302_219_fu_30362_p3;
wire   [31:0] select_ln350_109_fu_30370_p3;
wire  signed [31:0] lhs_92_fu_29572_p3;
wire  signed [31:0] rhs_110_fu_26033_p3;
wire  signed [32:0] sext_ln813_204_fu_30390_p1;
wire  signed [32:0] sext_ln813_203_fu_30386_p1;
wire   [32:0] ret_V_110_fu_30394_p2;
wire   [31:0] p_Val2_705_fu_30408_p2;
wire   [0:0] p_Result_705_fu_30400_p3;
wire   [0:0] p_Result_706_fu_30414_p3;
wire   [0:0] xor_ln895_434_fu_30422_p2;
wire   [0:0] xor_ln896_434_fu_30434_p2;
wire   [0:0] xor_ln302_221_fu_30446_p2;
wire   [0:0] overflow_272_fu_30428_p2;
wire   [0:0] xor_ln302_222_fu_30452_p2;
wire   [0:0] underflow_272_fu_30440_p2;
wire   [0:0] or_ln302_110_fu_30458_p2;
wire   [31:0] select_ln302_221_fu_30464_p3;
wire   [31:0] select_ln350_110_fu_30472_p3;
wire  signed [31:0] lhs_93_fu_29672_p3;
wire  signed [31:0] rhs_111_fu_26158_p3;
wire  signed [32:0] sext_ln813_206_fu_30492_p1;
wire  signed [32:0] sext_ln813_205_fu_30488_p1;
wire   [32:0] ret_V_111_fu_30496_p2;
wire   [31:0] p_Val2_707_fu_30510_p2;
wire   [0:0] p_Result_707_fu_30502_p3;
wire   [0:0] p_Result_708_fu_30516_p3;
wire   [0:0] xor_ln895_435_fu_30524_p2;
wire   [0:0] xor_ln896_435_fu_30536_p2;
wire   [0:0] xor_ln302_223_fu_30548_p2;
wire   [0:0] overflow_273_fu_30530_p2;
wire   [0:0] xor_ln302_224_fu_30554_p2;
wire   [0:0] underflow_273_fu_30542_p2;
wire   [0:0] or_ln302_111_fu_30560_p2;
wire   [31:0] select_ln302_223_fu_30566_p3;
wire   [31:0] select_ln350_111_fu_30574_p3;
wire  signed [31:0] lhs_94_fu_29772_p3;
wire  signed [31:0] rhs_112_fu_26283_p3;
wire  signed [32:0] sext_ln813_208_fu_30594_p1;
wire  signed [32:0] sext_ln813_207_fu_30590_p1;
wire   [32:0] ret_V_112_fu_30598_p2;
wire   [31:0] p_Val2_709_fu_30612_p2;
wire   [0:0] p_Result_709_fu_30604_p3;
wire   [0:0] p_Result_710_fu_30618_p3;
wire   [0:0] xor_ln895_436_fu_30626_p2;
wire   [0:0] xor_ln896_436_fu_30638_p2;
wire   [0:0] xor_ln302_225_fu_30650_p2;
wire   [0:0] overflow_274_fu_30632_p2;
wire   [0:0] xor_ln302_226_fu_30656_p2;
wire   [0:0] underflow_274_fu_30644_p2;
wire   [0:0] or_ln302_112_fu_30662_p2;
wire   [31:0] select_ln302_225_fu_30668_p3;
wire   [31:0] select_ln350_112_fu_30676_p3;
wire  signed [31:0] lhs_95_fu_29872_p3;
wire  signed [31:0] rhs_113_fu_26301_p3;
wire  signed [32:0] sext_ln813_210_fu_30696_p1;
wire  signed [32:0] sext_ln813_209_fu_30692_p1;
wire   [32:0] ret_V_113_fu_30700_p2;
wire   [31:0] p_Val2_711_fu_30714_p2;
wire   [0:0] p_Result_711_fu_30706_p3;
wire   [0:0] p_Result_712_fu_30720_p3;
wire   [0:0] xor_ln895_437_fu_30728_p2;
wire   [0:0] xor_ln896_437_fu_30740_p2;
wire   [0:0] xor_ln302_227_fu_30752_p2;
wire   [0:0] overflow_275_fu_30734_p2;
wire   [0:0] xor_ln302_228_fu_30758_p2;
wire   [0:0] underflow_275_fu_30746_p2;
wire   [0:0] or_ln302_113_fu_30764_p2;
wire   [31:0] select_ln302_227_fu_30770_p3;
wire   [31:0] select_ln350_113_fu_30778_p3;
wire  signed [31:0] lhs_96_fu_29972_p3;
wire  signed [31:0] rhs_114_fu_26425_p3;
wire  signed [32:0] sext_ln813_212_fu_30798_p1;
wire  signed [32:0] sext_ln813_211_fu_30794_p1;
wire   [32:0] ret_V_114_fu_30802_p2;
wire   [31:0] p_Val2_713_fu_30816_p2;
wire   [0:0] p_Result_713_fu_30808_p3;
wire   [0:0] p_Result_714_fu_30822_p3;
wire   [0:0] xor_ln895_438_fu_30830_p2;
wire   [0:0] xor_ln896_438_fu_30842_p2;
wire   [0:0] xor_ln302_229_fu_30854_p2;
wire   [0:0] overflow_276_fu_30836_p2;
wire   [0:0] xor_ln302_230_fu_30860_p2;
wire   [0:0] underflow_276_fu_30848_p2;
wire   [0:0] or_ln302_114_fu_30866_p2;
wire   [31:0] select_ln302_229_fu_30872_p3;
wire   [31:0] select_ln350_114_fu_30880_p3;
wire  signed [31:0] lhs_97_fu_30072_p3;
wire  signed [31:0] rhs_115_fu_26550_p3;
wire  signed [32:0] sext_ln813_214_fu_30900_p1;
wire  signed [32:0] sext_ln813_213_fu_30896_p1;
wire   [32:0] ret_V_115_fu_30904_p2;
wire   [31:0] p_Val2_715_fu_30918_p2;
wire   [0:0] p_Result_715_fu_30910_p3;
wire   [0:0] p_Result_716_fu_30924_p3;
wire   [0:0] xor_ln895_439_fu_30932_p2;
wire   [0:0] xor_ln896_439_fu_30944_p2;
wire   [0:0] xor_ln302_231_fu_30956_p2;
wire   [0:0] overflow_277_fu_30938_p2;
wire   [0:0] xor_ln302_232_fu_30962_p2;
wire   [0:0] underflow_277_fu_30950_p2;
wire   [0:0] or_ln302_115_fu_30968_p2;
wire   [31:0] select_ln302_231_fu_30974_p3;
wire   [31:0] select_ln350_115_fu_30982_p3;
wire  signed [31:0] lhs_98_fu_30174_p3;
wire  signed [31:0] rhs_116_fu_26695_p3;
wire  signed [32:0] sext_ln813_216_fu_31002_p1;
wire  signed [32:0] sext_ln813_215_fu_30998_p1;
wire   [32:0] ret_V_116_fu_31006_p2;
wire  signed [31:0] lhs_99_fu_30276_p3;
wire  signed [31:0] rhs_117_fu_26844_p3;
wire  signed [32:0] sext_ln813_218_fu_31038_p1;
wire  signed [32:0] sext_ln813_217_fu_31034_p1;
wire   [32:0] ret_V_117_fu_31042_p2;
wire  signed [31:0] lhs_100_fu_30378_p3;
wire  signed [31:0] rhs_118_fu_26993_p3;
wire  signed [32:0] sext_ln813_220_fu_31074_p1;
wire  signed [32:0] sext_ln813_219_fu_31070_p1;
wire   [32:0] ret_V_118_fu_31078_p2;
wire  signed [31:0] lhs_101_fu_30480_p3;
wire  signed [31:0] rhs_119_fu_27142_p3;
wire  signed [32:0] sext_ln813_222_fu_31110_p1;
wire  signed [32:0] sext_ln813_221_fu_31106_p1;
wire   [32:0] ret_V_119_fu_31114_p2;
wire  signed [31:0] lhs_102_fu_30582_p3;
wire  signed [31:0] rhs_120_fu_27291_p3;
wire  signed [32:0] sext_ln813_224_fu_31146_p1;
wire  signed [32:0] sext_ln813_223_fu_31142_p1;
wire   [32:0] ret_V_120_fu_31150_p2;
wire  signed [31:0] lhs_103_fu_30684_p3;
wire  signed [31:0] rhs_121_fu_27440_p3;
wire  signed [32:0] sext_ln813_226_fu_31182_p1;
wire  signed [32:0] sext_ln813_225_fu_31178_p1;
wire   [32:0] ret_V_121_fu_31186_p2;
wire  signed [31:0] lhs_104_fu_30786_p3;
wire  signed [31:0] rhs_122_fu_27589_p3;
wire  signed [32:0] sext_ln813_228_fu_31218_p1;
wire  signed [32:0] sext_ln813_227_fu_31214_p1;
wire   [32:0] ret_V_122_fu_31222_p2;
wire  signed [31:0] lhs_105_fu_30888_p3;
wire  signed [31:0] rhs_123_fu_27738_p3;
wire  signed [32:0] sext_ln813_230_fu_31254_p1;
wire  signed [32:0] sext_ln813_229_fu_31250_p1;
wire   [32:0] ret_V_123_fu_31258_p2;
wire  signed [31:0] lhs_106_fu_30990_p3;
wire  signed [31:0] rhs_124_fu_27887_p3;
wire  signed [32:0] sext_ln813_232_fu_31290_p1;
wire  signed [32:0] sext_ln813_231_fu_31286_p1;
wire   [32:0] ret_V_124_fu_31294_p2;
wire   [31:0] select_ln346_207_fu_31325_p3;
wire  signed [31:0] sext_ln856_119_fu_31322_p1;
wire   [0:0] xor_ln896_334_fu_31342_p2;
wire   [0:0] xor_ln888_250_fu_31352_p2;
wire   [0:0] or_ln888_126_fu_31357_p2;
wire   [0:0] tmp_918_fu_31367_p3;
wire   [0:0] xor_ln890_124_fu_31375_p2;
wire   [0:0] or_ln890_126_fu_31381_p2;
wire   [0:0] carry_251_fu_31347_p2;
wire   [0:0] deleted_zeros_123_fu_31362_p2;
wire   [0:0] xor_ln895_334_fu_31397_p2;
wire   [0:0] or_ln895_126_fu_31403_p2;
wire   [0:0] xor_ln895_335_fu_31408_p2;
wire   [0:0] deleted_ones_207_fu_31387_p2;
wire   [0:0] xor_ln896_335_fu_31419_p2;
wire   [0:0] and_ln891_126_fu_31392_p2;
wire   [0:0] or_ln896_126_fu_31425_p2;
wire   [0:0] xor_ln896_531_fu_31431_p2;
wire   [0:0] overflow_207_fu_31413_p2;
wire   [0:0] underflow_207_fu_31437_p2;
wire   [0:0] or_ln346_126_fu_31450_p2;
wire   [31:0] select_ln346_208_fu_31442_p3;
wire  signed [31:0] sext_ln856_120_fu_31339_p1;
wire   [0:0] xor_ln896_336_fu_31467_p2;
wire   [0:0] xor_ln888_252_fu_31477_p2;
wire   [0:0] or_ln888_127_fu_31482_p2;
wire   [0:0] tmp_924_fu_31492_p3;
wire   [0:0] xor_ln890_125_fu_31500_p2;
wire   [0:0] or_ln890_127_fu_31506_p2;
wire   [0:0] carry_253_fu_31472_p2;
wire   [0:0] deleted_zeros_124_fu_31487_p2;
wire   [0:0] xor_ln895_336_fu_31522_p2;
wire   [0:0] or_ln895_127_fu_31528_p2;
wire   [0:0] xor_ln895_337_fu_31533_p2;
wire   [0:0] deleted_ones_208_fu_31512_p2;
wire   [0:0] xor_ln896_337_fu_31544_p2;
wire   [0:0] and_ln891_127_fu_31517_p2;
wire   [0:0] or_ln896_127_fu_31550_p2;
wire   [0:0] xor_ln896_532_fu_31556_p2;
wire   [0:0] overflow_208_fu_31538_p2;
wire   [0:0] underflow_208_fu_31562_p2;
wire   [0:0] or_ln346_127_fu_31575_p2;
wire   [31:0] select_ln346_209_fu_31567_p3;
wire  signed [31:0] sext_ln856_121_fu_31464_p1;
wire   [0:0] xor_ln896_338_fu_31592_p2;
wire   [0:0] xor_ln888_254_fu_31602_p2;
wire   [0:0] or_ln888_128_fu_31607_p2;
wire   [0:0] tmp_930_fu_31617_p3;
wire   [0:0] xor_ln890_126_fu_31625_p2;
wire   [0:0] or_ln890_128_fu_31631_p2;
wire   [0:0] carry_255_fu_31597_p2;
wire   [0:0] deleted_zeros_125_fu_31612_p2;
wire   [0:0] xor_ln895_338_fu_31647_p2;
wire   [0:0] or_ln895_128_fu_31653_p2;
wire   [0:0] xor_ln895_339_fu_31658_p2;
wire   [0:0] deleted_ones_209_fu_31637_p2;
wire   [0:0] xor_ln896_339_fu_31669_p2;
wire   [0:0] and_ln891_128_fu_31642_p2;
wire   [0:0] or_ln896_128_fu_31675_p2;
wire   [0:0] xor_ln896_533_fu_31681_p2;
wire   [0:0] overflow_209_fu_31663_p2;
wire   [0:0] underflow_209_fu_31687_p2;
wire   [0:0] or_ln346_128_fu_31700_p2;
wire   [31:0] select_ln346_210_fu_31692_p3;
wire  signed [31:0] sext_ln856_122_fu_31589_p1;
wire   [0:0] xor_ln896_340_fu_31717_p2;
wire   [0:0] xor_ln888_256_fu_31727_p2;
wire   [0:0] or_ln888_129_fu_31732_p2;
wire   [0:0] tmp_936_fu_31742_p3;
wire   [0:0] xor_ln890_127_fu_31750_p2;
wire   [0:0] or_ln890_129_fu_31756_p2;
wire   [0:0] carry_257_fu_31722_p2;
wire   [0:0] deleted_zeros_126_fu_31737_p2;
wire   [0:0] xor_ln895_340_fu_31772_p2;
wire   [0:0] or_ln895_129_fu_31778_p2;
wire   [0:0] xor_ln895_341_fu_31783_p2;
wire   [0:0] deleted_ones_210_fu_31762_p2;
wire   [0:0] xor_ln896_341_fu_31794_p2;
wire   [0:0] and_ln891_129_fu_31767_p2;
wire   [0:0] or_ln896_129_fu_31800_p2;
wire   [0:0] xor_ln896_534_fu_31806_p2;
wire   [0:0] overflow_210_fu_31788_p2;
wire   [0:0] underflow_210_fu_31812_p2;
wire   [0:0] or_ln346_129_fu_31825_p2;
wire   [31:0] select_ln346_211_fu_31817_p3;
wire  signed [31:0] sext_ln856_123_fu_31714_p1;
wire   [0:0] xor_ln896_342_fu_31842_p2;
wire   [0:0] xor_ln888_258_fu_31852_p2;
wire   [0:0] or_ln888_130_fu_31857_p2;
wire   [0:0] tmp_942_fu_31867_p3;
wire   [0:0] xor_ln890_128_fu_31875_p2;
wire   [0:0] or_ln890_130_fu_31881_p2;
wire   [0:0] carry_259_fu_31847_p2;
wire   [0:0] deleted_zeros_127_fu_31862_p2;
wire   [0:0] xor_ln895_342_fu_31897_p2;
wire   [0:0] or_ln895_130_fu_31903_p2;
wire   [0:0] xor_ln895_343_fu_31908_p2;
wire   [0:0] deleted_ones_211_fu_31887_p2;
wire   [0:0] xor_ln896_343_fu_31919_p2;
wire   [0:0] and_ln891_130_fu_31892_p2;
wire   [0:0] or_ln896_130_fu_31925_p2;
wire   [0:0] xor_ln896_535_fu_31931_p2;
wire   [0:0] overflow_211_fu_31913_p2;
wire   [0:0] underflow_211_fu_31937_p2;
wire   [0:0] or_ln346_130_fu_31950_p2;
wire   [31:0] select_ln346_212_fu_31942_p3;
wire  signed [31:0] sext_ln856_124_fu_31839_p1;
wire   [0:0] xor_ln896_344_fu_31967_p2;
wire   [0:0] xor_ln888_260_fu_31977_p2;
wire   [0:0] or_ln888_131_fu_31982_p2;
wire   [0:0] tmp_948_fu_31992_p3;
wire   [0:0] xor_ln890_129_fu_32000_p2;
wire   [0:0] or_ln890_131_fu_32006_p2;
wire   [0:0] carry_261_fu_31972_p2;
wire   [0:0] deleted_zeros_128_fu_31987_p2;
wire   [0:0] xor_ln895_344_fu_32022_p2;
wire   [0:0] or_ln895_131_fu_32028_p2;
wire   [0:0] xor_ln895_345_fu_32033_p2;
wire   [0:0] deleted_ones_212_fu_32012_p2;
wire   [0:0] xor_ln896_345_fu_32044_p2;
wire   [0:0] and_ln891_131_fu_32017_p2;
wire   [0:0] or_ln896_131_fu_32050_p2;
wire   [0:0] xor_ln896_536_fu_32056_p2;
wire   [0:0] overflow_212_fu_32038_p2;
wire   [0:0] underflow_212_fu_32062_p2;
wire   [0:0] or_ln346_131_fu_32075_p2;
wire   [31:0] select_ln346_213_fu_32067_p3;
wire  signed [31:0] sext_ln856_125_fu_31964_p1;
wire   [0:0] xor_ln896_346_fu_32092_p2;
wire   [0:0] xor_ln888_262_fu_32102_p2;
wire   [0:0] or_ln888_132_fu_32107_p2;
wire   [0:0] tmp_954_fu_32117_p3;
wire   [0:0] xor_ln890_130_fu_32125_p2;
wire   [0:0] or_ln890_132_fu_32131_p2;
wire   [0:0] carry_263_fu_32097_p2;
wire   [0:0] deleted_zeros_129_fu_32112_p2;
wire   [0:0] xor_ln895_346_fu_32147_p2;
wire   [0:0] or_ln895_132_fu_32153_p2;
wire   [0:0] xor_ln895_347_fu_32158_p2;
wire   [0:0] deleted_ones_213_fu_32137_p2;
wire   [0:0] xor_ln896_347_fu_32169_p2;
wire   [0:0] and_ln891_132_fu_32142_p2;
wire   [0:0] or_ln896_132_fu_32175_p2;
wire   [0:0] xor_ln896_537_fu_32181_p2;
wire   [0:0] overflow_213_fu_32163_p2;
wire   [0:0] underflow_213_fu_32187_p2;
wire   [0:0] or_ln346_132_fu_32200_p2;
wire   [31:0] select_ln346_214_fu_32192_p3;
wire  signed [31:0] sext_ln856_126_fu_32089_p1;
wire   [0:0] xor_ln896_348_fu_32217_p2;
wire   [0:0] xor_ln888_264_fu_32227_p2;
wire   [0:0] or_ln888_133_fu_32232_p2;
wire   [0:0] tmp_960_fu_32242_p3;
wire   [0:0] xor_ln890_131_fu_32250_p2;
wire   [0:0] or_ln890_133_fu_32256_p2;
wire   [0:0] carry_265_fu_32222_p2;
wire   [0:0] deleted_zeros_130_fu_32237_p2;
wire   [0:0] xor_ln895_348_fu_32272_p2;
wire   [0:0] or_ln895_133_fu_32278_p2;
wire   [0:0] xor_ln895_349_fu_32283_p2;
wire   [0:0] deleted_ones_214_fu_32262_p2;
wire   [0:0] xor_ln896_349_fu_32294_p2;
wire   [0:0] and_ln891_133_fu_32267_p2;
wire   [0:0] or_ln896_133_fu_32300_p2;
wire   [0:0] xor_ln896_538_fu_32306_p2;
wire   [0:0] overflow_214_fu_32288_p2;
wire   [0:0] underflow_214_fu_32312_p2;
wire   [0:0] or_ln346_133_fu_32325_p2;
wire   [31:0] select_ln346_215_fu_32317_p3;
wire  signed [31:0] sext_ln856_127_fu_32214_p1;
wire   [20:0] zext_ln377_134_fu_32342_p1;
wire  signed [20:0] sext_ln823_128_fu_32339_p1;
wire  signed [20:0] p_Val2_565_fu_32345_p2;
wire   [0:0] p_Result_566_fu_32355_p3;
wire   [0:0] xor_ln896_350_fu_32363_p2;
wire   [0:0] xor_ln888_266_fu_32374_p2;
wire   [0:0] or_ln888_134_fu_32379_p2;
wire   [0:0] tmp_966_fu_32390_p3;
wire   [0:0] xor_ln890_132_fu_32398_p2;
wire   [0:0] or_ln890_134_fu_32404_p2;
wire   [0:0] carry_267_fu_32369_p2;
wire   [0:0] deleted_zeros_131_fu_32385_p2;
wire   [0:0] xor_ln895_350_fu_32420_p2;
wire   [0:0] or_ln895_134_fu_32426_p2;
wire   [0:0] xor_ln895_351_fu_32432_p2;
wire   [0:0] deleted_ones_215_fu_32410_p2;
wire   [0:0] xor_ln896_351_fu_32443_p2;
wire   [0:0] and_ln891_134_fu_32415_p2;
wire   [0:0] or_ln896_134_fu_32449_p2;
wire   [0:0] xor_ln896_539_fu_32455_p2;
wire   [0:0] overflow_215_fu_32437_p2;
wire   [0:0] underflow_215_fu_32461_p2;
wire   [0:0] or_ln346_134_fu_32474_p2;
wire   [31:0] select_ln346_216_fu_32466_p3;
wire  signed [31:0] sext_ln856_128_fu_32351_p1;
wire   [19:0] zext_ln377_135_fu_32491_p1;
wire  signed [19:0] sext_ln823_129_fu_32488_p1;
wire  signed [19:0] p_Val2_568_fu_32494_p2;
wire   [0:0] p_Result_569_fu_32504_p3;
wire   [0:0] xor_ln896_352_fu_32512_p2;
wire   [0:0] xor_ln888_268_fu_32523_p2;
wire   [0:0] or_ln888_135_fu_32528_p2;
wire   [0:0] tmp_972_fu_32539_p3;
wire   [0:0] xor_ln890_133_fu_32547_p2;
wire   [0:0] or_ln890_135_fu_32553_p2;
wire   [0:0] carry_269_fu_32518_p2;
wire   [0:0] deleted_zeros_132_fu_32534_p2;
wire   [0:0] xor_ln895_352_fu_32569_p2;
wire   [0:0] or_ln895_135_fu_32575_p2;
wire   [0:0] xor_ln895_353_fu_32581_p2;
wire   [0:0] deleted_ones_216_fu_32559_p2;
wire   [0:0] xor_ln896_353_fu_32592_p2;
wire   [0:0] and_ln891_135_fu_32564_p2;
wire   [0:0] or_ln896_135_fu_32598_p2;
wire   [0:0] xor_ln896_540_fu_32604_p2;
wire   [0:0] overflow_216_fu_32586_p2;
wire   [0:0] underflow_216_fu_32610_p2;
wire   [0:0] or_ln346_135_fu_32623_p2;
wire   [31:0] select_ln346_217_fu_32615_p3;
wire  signed [31:0] sext_ln856_129_fu_32500_p1;
wire   [19:0] zext_ln377_136_fu_32640_p1;
wire  signed [19:0] sext_ln823_130_fu_32637_p1;
wire  signed [19:0] p_Val2_571_fu_32643_p2;
wire   [0:0] p_Result_572_fu_32653_p3;
wire   [0:0] xor_ln896_354_fu_32661_p2;
wire   [0:0] xor_ln888_270_fu_32672_p2;
wire   [0:0] or_ln888_136_fu_32677_p2;
wire   [0:0] tmp_978_fu_32688_p3;
wire   [0:0] xor_ln890_134_fu_32696_p2;
wire   [0:0] or_ln890_136_fu_32702_p2;
wire   [0:0] carry_271_fu_32667_p2;
wire   [0:0] deleted_zeros_133_fu_32683_p2;
wire   [0:0] xor_ln895_354_fu_32718_p2;
wire   [0:0] or_ln895_136_fu_32724_p2;
wire   [0:0] xor_ln895_355_fu_32730_p2;
wire   [0:0] deleted_ones_217_fu_32708_p2;
wire   [0:0] xor_ln896_355_fu_32741_p2;
wire   [0:0] and_ln891_136_fu_32713_p2;
wire   [0:0] or_ln896_136_fu_32747_p2;
wire   [0:0] xor_ln896_541_fu_32753_p2;
wire   [0:0] overflow_217_fu_32735_p2;
wire   [0:0] underflow_217_fu_32759_p2;
wire   [0:0] or_ln346_136_fu_32772_p2;
wire   [31:0] select_ln346_218_fu_32764_p3;
wire  signed [31:0] sext_ln856_130_fu_32649_p1;
wire   [20:0] zext_ln377_137_fu_32789_p1;
wire  signed [20:0] sext_ln823_131_fu_32786_p1;
wire  signed [20:0] p_Val2_574_fu_32792_p2;
wire   [0:0] p_Result_575_fu_32802_p3;
wire   [0:0] xor_ln896_356_fu_32810_p2;
wire   [0:0] xor_ln888_272_fu_32821_p2;
wire   [0:0] or_ln888_137_fu_32826_p2;
wire   [0:0] tmp_984_fu_32837_p3;
wire   [0:0] xor_ln890_135_fu_32845_p2;
wire   [0:0] or_ln890_137_fu_32851_p2;
wire   [0:0] carry_273_fu_32816_p2;
wire   [0:0] deleted_zeros_134_fu_32832_p2;
wire   [0:0] xor_ln895_356_fu_32867_p2;
wire   [0:0] or_ln895_137_fu_32873_p2;
wire   [0:0] xor_ln895_357_fu_32879_p2;
wire   [0:0] deleted_ones_218_fu_32857_p2;
wire   [0:0] xor_ln896_357_fu_32890_p2;
wire   [0:0] and_ln891_137_fu_32862_p2;
wire   [0:0] or_ln896_137_fu_32896_p2;
wire   [0:0] xor_ln896_542_fu_32902_p2;
wire   [0:0] overflow_218_fu_32884_p2;
wire   [0:0] underflow_218_fu_32908_p2;
wire   [0:0] or_ln346_137_fu_32921_p2;
wire   [31:0] select_ln346_219_fu_32913_p3;
wire  signed [31:0] sext_ln856_131_fu_32798_p1;
wire   [19:0] zext_ln377_138_fu_32938_p1;
wire  signed [19:0] sext_ln823_132_fu_32935_p1;
wire  signed [19:0] p_Val2_577_fu_32941_p2;
wire   [0:0] p_Result_578_fu_32951_p3;
wire   [0:0] xor_ln896_358_fu_32959_p2;
wire   [0:0] xor_ln888_274_fu_32970_p2;
wire   [0:0] or_ln888_138_fu_32975_p2;
wire   [0:0] tmp_990_fu_32986_p3;
wire   [0:0] xor_ln890_136_fu_32994_p2;
wire   [0:0] or_ln890_138_fu_33000_p2;
wire   [0:0] carry_275_fu_32965_p2;
wire   [0:0] deleted_zeros_135_fu_32981_p2;
wire   [0:0] xor_ln895_358_fu_33016_p2;
wire   [0:0] or_ln895_138_fu_33022_p2;
wire   [0:0] xor_ln895_359_fu_33028_p2;
wire   [0:0] deleted_ones_219_fu_33006_p2;
wire   [0:0] xor_ln896_359_fu_33039_p2;
wire   [0:0] and_ln891_138_fu_33011_p2;
wire   [0:0] or_ln896_138_fu_33045_p2;
wire   [0:0] xor_ln896_543_fu_33051_p2;
wire   [0:0] overflow_219_fu_33033_p2;
wire   [0:0] underflow_219_fu_33057_p2;
wire   [0:0] or_ln346_138_fu_33070_p2;
wire   [31:0] select_ln346_220_fu_33062_p3;
wire  signed [31:0] sext_ln856_132_fu_32947_p1;
wire   [19:0] zext_ln377_139_fu_33087_p1;
wire  signed [19:0] sext_ln823_133_fu_33084_p1;
wire  signed [19:0] p_Val2_580_fu_33090_p2;
wire   [0:0] p_Result_581_fu_33100_p3;
wire   [0:0] xor_ln896_360_fu_33108_p2;
wire   [0:0] xor_ln888_276_fu_33119_p2;
wire   [0:0] or_ln888_139_fu_33124_p2;
wire   [0:0] tmp_996_fu_33135_p3;
wire   [0:0] xor_ln890_137_fu_33143_p2;
wire   [0:0] or_ln890_139_fu_33149_p2;
wire   [0:0] carry_277_fu_33114_p2;
wire   [0:0] deleted_zeros_136_fu_33130_p2;
wire   [0:0] xor_ln895_360_fu_33165_p2;
wire   [0:0] or_ln895_139_fu_33171_p2;
wire   [0:0] xor_ln895_361_fu_33177_p2;
wire   [0:0] deleted_ones_220_fu_33155_p2;
wire   [0:0] xor_ln896_361_fu_33188_p2;
wire   [0:0] and_ln891_139_fu_33160_p2;
wire   [0:0] or_ln896_139_fu_33194_p2;
wire   [0:0] xor_ln896_544_fu_33200_p2;
wire   [0:0] overflow_220_fu_33182_p2;
wire   [0:0] underflow_220_fu_33206_p2;
wire   [0:0] or_ln346_139_fu_33219_p2;
wire   [31:0] select_ln346_221_fu_33211_p3;
wire  signed [31:0] sext_ln856_133_fu_33096_p1;
wire   [17:0] zext_ln377_140_fu_33236_p1;
wire  signed [17:0] sext_ln823_134_fu_33233_p1;
wire  signed [17:0] p_Val2_583_fu_33239_p2;
wire   [0:0] p_Result_584_fu_33249_p3;
wire   [0:0] xor_ln896_362_fu_33257_p2;
wire   [0:0] xor_ln888_278_fu_33268_p2;
wire   [0:0] or_ln888_140_fu_33273_p2;
wire   [0:0] tmp_1002_fu_33284_p3;
wire   [0:0] xor_ln890_138_fu_33292_p2;
wire   [0:0] or_ln890_140_fu_33298_p2;
wire   [0:0] carry_279_fu_33263_p2;
wire   [0:0] deleted_zeros_137_fu_33279_p2;
wire   [0:0] xor_ln895_362_fu_33314_p2;
wire   [0:0] or_ln895_140_fu_33320_p2;
wire   [0:0] xor_ln895_363_fu_33326_p2;
wire   [0:0] deleted_ones_221_fu_33304_p2;
wire   [0:0] xor_ln896_363_fu_33337_p2;
wire   [0:0] and_ln891_140_fu_33309_p2;
wire   [0:0] or_ln896_140_fu_33343_p2;
wire   [0:0] xor_ln896_545_fu_33349_p2;
wire   [0:0] overflow_221_fu_33331_p2;
wire   [0:0] underflow_221_fu_33355_p2;
wire   [0:0] or_ln346_140_fu_33368_p2;
wire   [31:0] select_ln346_222_fu_33360_p3;
wire  signed [31:0] sext_ln856_134_fu_33245_p1;
wire   [18:0] zext_ln377_141_fu_33385_p1;
wire  signed [18:0] sext_ln823_135_fu_33382_p1;
wire  signed [18:0] p_Val2_586_fu_33388_p2;
wire   [0:0] p_Result_587_fu_33398_p3;
wire   [0:0] xor_ln896_364_fu_33406_p2;
wire   [0:0] xor_ln888_280_fu_33417_p2;
wire   [0:0] or_ln888_141_fu_33422_p2;
wire   [0:0] tmp_1008_fu_33433_p3;
wire   [0:0] xor_ln890_139_fu_33441_p2;
wire   [0:0] or_ln890_141_fu_33447_p2;
wire   [0:0] carry_281_fu_33412_p2;
wire   [0:0] deleted_zeros_138_fu_33428_p2;
wire   [0:0] xor_ln895_364_fu_33463_p2;
wire   [0:0] or_ln895_141_fu_33469_p2;
wire   [0:0] xor_ln895_365_fu_33475_p2;
wire   [0:0] deleted_ones_222_fu_33453_p2;
wire   [0:0] xor_ln896_365_fu_33486_p2;
wire   [0:0] and_ln891_141_fu_33458_p2;
wire   [0:0] or_ln896_141_fu_33492_p2;
wire   [0:0] xor_ln896_546_fu_33498_p2;
wire   [0:0] overflow_222_fu_33480_p2;
wire   [0:0] underflow_222_fu_33504_p2;
wire   [0:0] or_ln346_141_fu_33517_p2;
wire   [31:0] select_ln346_223_fu_33509_p3;
wire  signed [31:0] sext_ln856_135_fu_33394_p1;
wire   [31:0] select_ln346_224_fu_33534_p3;
wire  signed [31:0] sext_ln856_136_fu_33531_p1;
wire   [30:0] p_Val2_591_fu_33580_p4;
wire   [0:0] tmp_1017_fu_33602_p3;
wire   [31:0] zext_ln377_143_fu_33610_p1;
wire  signed [31:0] sext_ln818_2_fu_33590_p1;
wire   [19:0] p_Val2_594_fu_33644_p4;
wire   [0:0] tmp_1023_fu_33666_p3;
wire   [20:0] zext_ln377_144_fu_33674_p1;
wire  signed [20:0] sext_ln823_137_fu_33654_p1;
wire   [18:0] p_Val2_597_fu_33708_p4;
wire   [0:0] tmp_1029_fu_33730_p3;
wire   [19:0] zext_ln377_145_fu_33738_p1;
wire  signed [19:0] sext_ln823_138_fu_33718_p1;
wire   [25:0] p_Val2_600_fu_33772_p4;
wire   [0:0] tmp_1035_fu_33794_p3;
wire   [26:0] zext_ln377_146_fu_33802_p1;
wire  signed [26:0] sext_ln823_139_fu_33782_p1;
wire   [24:0] p_Val2_603_fu_33836_p4;
wire   [0:0] tmp_1041_fu_33858_p3;
wire   [25:0] zext_ln377_147_fu_33866_p1;
wire  signed [25:0] sext_ln823_140_fu_33846_p1;
wire   [19:0] p_Val2_606_fu_33900_p4;
wire   [0:0] tmp_1047_fu_33922_p3;
wire   [20:0] zext_ln377_148_fu_33930_p1;
wire  signed [20:0] sext_ln823_141_fu_33910_p1;
wire   [19:0] p_Val2_609_fu_33964_p4;
wire   [0:0] tmp_1053_fu_33986_p3;
wire   [20:0] zext_ln377_149_fu_33994_p1;
wire  signed [20:0] sext_ln823_142_fu_33974_p1;
wire   [19:0] p_Val2_612_fu_34028_p4;
wire   [0:0] tmp_1059_fu_34050_p3;
wire   [20:0] zext_ln377_150_fu_34058_p1;
wire  signed [20:0] sext_ln823_143_fu_34038_p1;
wire   [24:0] p_Val2_615_fu_34092_p4;
wire   [0:0] tmp_1065_fu_34114_p3;
wire   [25:0] zext_ln377_151_fu_34122_p1;
wire  signed [25:0] sext_ln823_144_fu_34102_p1;
wire   [34:0] shl_ln1273_18_fu_34462_p3;
wire  signed [35:0] sext_ln1273_20_fu_34469_p1;
wire   [32:0] shl_ln1273_19_fu_34479_p3;
wire   [35:0] sub_ln1273_10_fu_34473_p2;
wire  signed [35:0] sext_ln1273_21_fu_34486_p1;
wire   [35:0] r_V_156_fu_34490_p2;
wire   [11:0] p_Val2_639_fu_34504_p4;
wire   [0:0] tmp_1113_fu_34526_p3;
wire   [12:0] zext_ln377_159_fu_34534_p1;
wire  signed [12:0] sext_ln823_151_fu_34514_p1;
wire   [0:0] p_Result_641_fu_34544_p3;
wire   [0:0] p_Result_640_fu_34518_p3;
wire   [0:0] xor_ln896_400_fu_34552_p2;
wire   [0:0] xor_ln888_316_fu_34572_p2;
wire   [0:0] Range2_all_ones_157_fu_34564_p3;
wire   [0:0] or_ln888_159_fu_34578_p2;
wire   [0:0] tmp_1116_fu_34590_p3;
wire   [0:0] xor_ln890_157_fu_34598_p2;
wire   [0:0] or_ln890_159_fu_34604_p2;
wire   [0:0] carry_317_fu_34558_p2;
wire   [0:0] deleted_zeros_156_fu_34584_p2;
wire   [0:0] xor_ln895_400_fu_34622_p2;
wire   [0:0] p_Result_639_fu_34496_p3;
wire   [0:0] or_ln895_159_fu_34628_p2;
wire   [0:0] xor_ln895_401_fu_34634_p2;
wire   [0:0] deleted_ones_240_fu_34610_p2;
wire   [0:0] xor_ln896_401_fu_34646_p2;
wire   [0:0] and_ln891_159_fu_34616_p2;
wire   [0:0] or_ln896_159_fu_34652_p2;
wire   [0:0] xor_ln896_564_fu_34658_p2;
wire   [0:0] underflow_240_fu_34664_p2;
wire   [0:0] xor_ln895_440_fu_34718_p2;
wire   [0:0] xor_ln896_440_fu_34728_p2;
wire   [0:0] xor_ln302_233_fu_34738_p2;
wire   [0:0] overflow_278_fu_34723_p2;
wire   [0:0] xor_ln302_234_fu_34742_p2;
wire   [0:0] underflow_278_fu_34733_p2;
wire   [0:0] or_ln302_116_fu_34748_p2;
wire   [31:0] select_ln302_233_fu_34754_p3;
wire   [31:0] select_ln350_116_fu_34761_p3;
wire   [0:0] xor_ln895_441_fu_34776_p2;
wire   [0:0] xor_ln896_441_fu_34786_p2;
wire   [0:0] xor_ln302_235_fu_34796_p2;
wire   [0:0] overflow_279_fu_34781_p2;
wire   [0:0] xor_ln302_236_fu_34800_p2;
wire   [0:0] underflow_279_fu_34791_p2;
wire   [0:0] or_ln302_117_fu_34806_p2;
wire   [31:0] select_ln302_235_fu_34812_p3;
wire   [31:0] select_ln350_117_fu_34819_p3;
wire   [0:0] xor_ln895_442_fu_34834_p2;
wire   [0:0] xor_ln896_442_fu_34844_p2;
wire   [0:0] xor_ln302_237_fu_34854_p2;
wire   [0:0] overflow_280_fu_34839_p2;
wire   [0:0] xor_ln302_238_fu_34858_p2;
wire   [0:0] underflow_280_fu_34849_p2;
wire   [0:0] or_ln302_118_fu_34864_p2;
wire   [31:0] select_ln302_237_fu_34870_p3;
wire   [31:0] select_ln350_118_fu_34877_p3;
wire   [0:0] xor_ln895_443_fu_34892_p2;
wire   [0:0] xor_ln896_443_fu_34902_p2;
wire   [0:0] xor_ln302_239_fu_34912_p2;
wire   [0:0] overflow_281_fu_34897_p2;
wire   [0:0] xor_ln302_240_fu_34916_p2;
wire   [0:0] underflow_281_fu_34907_p2;
wire   [0:0] or_ln302_119_fu_34922_p2;
wire   [31:0] select_ln302_239_fu_34928_p3;
wire   [31:0] select_ln350_119_fu_34935_p3;
wire   [0:0] xor_ln895_444_fu_34950_p2;
wire   [0:0] xor_ln896_444_fu_34960_p2;
wire   [0:0] xor_ln302_241_fu_34970_p2;
wire   [0:0] overflow_282_fu_34955_p2;
wire   [0:0] xor_ln302_242_fu_34974_p2;
wire   [0:0] underflow_282_fu_34965_p2;
wire   [0:0] or_ln302_120_fu_34980_p2;
wire   [31:0] select_ln302_241_fu_34986_p3;
wire   [31:0] select_ln350_120_fu_34993_p3;
wire   [0:0] xor_ln895_445_fu_35008_p2;
wire   [0:0] xor_ln896_445_fu_35018_p2;
wire   [0:0] xor_ln302_243_fu_35028_p2;
wire   [0:0] overflow_283_fu_35013_p2;
wire   [0:0] xor_ln302_244_fu_35032_p2;
wire   [0:0] underflow_283_fu_35023_p2;
wire   [0:0] or_ln302_121_fu_35038_p2;
wire   [31:0] select_ln302_243_fu_35044_p3;
wire   [31:0] select_ln350_121_fu_35051_p3;
wire   [0:0] xor_ln895_446_fu_35066_p2;
wire   [0:0] xor_ln896_446_fu_35076_p2;
wire   [0:0] xor_ln302_245_fu_35086_p2;
wire   [0:0] overflow_284_fu_35071_p2;
wire   [0:0] xor_ln302_246_fu_35090_p2;
wire   [0:0] underflow_284_fu_35081_p2;
wire   [0:0] or_ln302_122_fu_35096_p2;
wire   [31:0] select_ln302_245_fu_35102_p3;
wire   [31:0] select_ln350_122_fu_35109_p3;
wire   [0:0] xor_ln895_447_fu_35124_p2;
wire   [0:0] xor_ln896_447_fu_35134_p2;
wire   [0:0] xor_ln302_247_fu_35144_p2;
wire   [0:0] overflow_285_fu_35129_p2;
wire   [0:0] xor_ln302_248_fu_35148_p2;
wire   [0:0] underflow_285_fu_35139_p2;
wire   [0:0] or_ln302_123_fu_35154_p2;
wire   [31:0] select_ln302_247_fu_35160_p3;
wire   [31:0] select_ln350_123_fu_35167_p3;
wire   [0:0] xor_ln895_448_fu_35182_p2;
wire   [0:0] xor_ln896_448_fu_35192_p2;
wire   [0:0] xor_ln302_249_fu_35202_p2;
wire   [0:0] overflow_286_fu_35187_p2;
wire   [0:0] xor_ln302_250_fu_35206_p2;
wire   [0:0] underflow_286_fu_35197_p2;
wire   [0:0] or_ln302_124_fu_35212_p2;
wire   [31:0] select_ln302_249_fu_35218_p3;
wire   [31:0] select_ln350_124_fu_35225_p3;
wire  signed [31:0] lhs_107_fu_34768_p3;
wire  signed [31:0] rhs_125_fu_31332_p3;
wire  signed [32:0] sext_ln813_234_fu_35244_p1;
wire  signed [32:0] sext_ln813_233_fu_35240_p1;
wire   [32:0] ret_V_125_fu_35248_p2;
wire   [31:0] p_Val2_735_fu_35262_p2;
wire   [0:0] p_Result_735_fu_35254_p3;
wire   [0:0] p_Result_736_fu_35268_p3;
wire   [0:0] xor_ln895_449_fu_35276_p2;
wire   [0:0] xor_ln896_449_fu_35288_p2;
wire   [0:0] xor_ln302_251_fu_35300_p2;
wire   [0:0] overflow_287_fu_35282_p2;
wire   [0:0] xor_ln302_252_fu_35306_p2;
wire   [0:0] underflow_287_fu_35294_p2;
wire   [0:0] or_ln302_125_fu_35312_p2;
wire   [31:0] select_ln302_251_fu_35318_p3;
wire   [31:0] select_ln350_125_fu_35326_p3;
wire  signed [31:0] lhs_108_fu_34826_p3;
wire  signed [31:0] rhs_126_fu_31456_p3;
wire  signed [32:0] sext_ln813_236_fu_35346_p1;
wire  signed [32:0] sext_ln813_235_fu_35342_p1;
wire   [32:0] ret_V_126_fu_35350_p2;
wire   [31:0] p_Val2_737_fu_35364_p2;
wire   [0:0] p_Result_737_fu_35356_p3;
wire   [0:0] p_Result_738_fu_35370_p3;
wire   [0:0] xor_ln895_450_fu_35378_p2;
wire   [0:0] xor_ln896_450_fu_35390_p2;
wire   [0:0] xor_ln302_253_fu_35402_p2;
wire   [0:0] overflow_288_fu_35384_p2;
wire   [0:0] xor_ln302_254_fu_35408_p2;
wire   [0:0] underflow_288_fu_35396_p2;
wire   [0:0] or_ln302_126_fu_35414_p2;
wire   [31:0] select_ln302_253_fu_35420_p3;
wire   [31:0] select_ln350_126_fu_35428_p3;
wire  signed [31:0] lhs_109_fu_34884_p3;
wire  signed [31:0] rhs_127_fu_31581_p3;
wire  signed [32:0] sext_ln813_238_fu_35448_p1;
wire  signed [32:0] sext_ln813_237_fu_35444_p1;
wire   [32:0] ret_V_127_fu_35452_p2;
wire   [31:0] p_Val2_739_fu_35466_p2;
wire   [0:0] p_Result_739_fu_35458_p3;
wire   [0:0] p_Result_740_fu_35472_p3;
wire   [0:0] xor_ln895_451_fu_35480_p2;
wire   [0:0] xor_ln896_451_fu_35492_p2;
wire   [0:0] xor_ln302_255_fu_35504_p2;
wire   [0:0] overflow_289_fu_35486_p2;
wire   [0:0] xor_ln302_256_fu_35510_p2;
wire   [0:0] underflow_289_fu_35498_p2;
wire   [0:0] or_ln302_127_fu_35516_p2;
wire   [31:0] select_ln302_255_fu_35522_p3;
wire   [31:0] select_ln350_127_fu_35530_p3;
wire  signed [31:0] lhs_110_fu_34942_p3;
wire  signed [31:0] rhs_128_fu_31706_p3;
wire  signed [32:0] sext_ln813_240_fu_35550_p1;
wire  signed [32:0] sext_ln813_239_fu_35546_p1;
wire   [32:0] ret_V_128_fu_35554_p2;
wire   [31:0] p_Val2_741_fu_35568_p2;
wire   [0:0] p_Result_741_fu_35560_p3;
wire   [0:0] p_Result_742_fu_35574_p3;
wire   [0:0] xor_ln895_452_fu_35582_p2;
wire   [0:0] xor_ln896_452_fu_35594_p2;
wire   [0:0] xor_ln302_257_fu_35606_p2;
wire   [0:0] overflow_290_fu_35588_p2;
wire   [0:0] xor_ln302_258_fu_35612_p2;
wire   [0:0] underflow_290_fu_35600_p2;
wire   [0:0] or_ln302_128_fu_35618_p2;
wire   [31:0] select_ln302_257_fu_35624_p3;
wire   [31:0] select_ln350_128_fu_35632_p3;
wire  signed [31:0] lhs_111_fu_35000_p3;
wire  signed [31:0] rhs_129_fu_31831_p3;
wire  signed [32:0] sext_ln813_242_fu_35652_p1;
wire  signed [32:0] sext_ln813_241_fu_35648_p1;
wire   [32:0] ret_V_129_fu_35656_p2;
wire   [31:0] p_Val2_743_fu_35670_p2;
wire   [0:0] p_Result_743_fu_35662_p3;
wire   [0:0] p_Result_744_fu_35676_p3;
wire   [0:0] xor_ln895_453_fu_35684_p2;
wire   [0:0] xor_ln896_453_fu_35696_p2;
wire   [0:0] xor_ln302_259_fu_35708_p2;
wire   [0:0] overflow_291_fu_35690_p2;
wire   [0:0] xor_ln302_260_fu_35714_p2;
wire   [0:0] underflow_291_fu_35702_p2;
wire   [0:0] or_ln302_129_fu_35720_p2;
wire   [31:0] select_ln302_259_fu_35726_p3;
wire   [31:0] select_ln350_129_fu_35734_p3;
wire  signed [31:0] lhs_112_fu_35058_p3;
wire  signed [31:0] rhs_130_fu_31956_p3;
wire  signed [32:0] sext_ln813_244_fu_35754_p1;
wire  signed [32:0] sext_ln813_243_fu_35750_p1;
wire   [32:0] ret_V_130_fu_35758_p2;
wire   [31:0] p_Val2_745_fu_35772_p2;
wire   [0:0] p_Result_745_fu_35764_p3;
wire   [0:0] p_Result_746_fu_35778_p3;
wire   [0:0] xor_ln895_454_fu_35786_p2;
wire   [0:0] xor_ln896_454_fu_35798_p2;
wire   [0:0] xor_ln302_261_fu_35810_p2;
wire   [0:0] overflow_292_fu_35792_p2;
wire   [0:0] xor_ln302_262_fu_35816_p2;
wire   [0:0] underflow_292_fu_35804_p2;
wire   [0:0] or_ln302_130_fu_35822_p2;
wire   [31:0] select_ln302_261_fu_35828_p3;
wire   [31:0] select_ln350_130_fu_35836_p3;
wire  signed [31:0] lhs_113_fu_35116_p3;
wire  signed [31:0] rhs_131_fu_32081_p3;
wire  signed [32:0] sext_ln813_246_fu_35856_p1;
wire  signed [32:0] sext_ln813_245_fu_35852_p1;
wire   [32:0] ret_V_131_fu_35860_p2;
wire   [31:0] p_Val2_747_fu_35874_p2;
wire   [0:0] p_Result_747_fu_35866_p3;
wire   [0:0] p_Result_748_fu_35880_p3;
wire   [0:0] xor_ln895_455_fu_35888_p2;
wire   [0:0] xor_ln896_455_fu_35900_p2;
wire   [0:0] xor_ln302_263_fu_35912_p2;
wire   [0:0] overflow_293_fu_35894_p2;
wire   [0:0] xor_ln302_264_fu_35918_p2;
wire   [0:0] underflow_293_fu_35906_p2;
wire   [0:0] or_ln302_131_fu_35924_p2;
wire   [31:0] select_ln302_263_fu_35930_p3;
wire   [31:0] select_ln350_131_fu_35938_p3;
wire  signed [31:0] lhs_114_fu_35174_p3;
wire  signed [31:0] rhs_132_fu_32206_p3;
wire  signed [32:0] sext_ln813_248_fu_35958_p1;
wire  signed [32:0] sext_ln813_247_fu_35954_p1;
wire   [32:0] ret_V_132_fu_35962_p2;
wire   [31:0] p_Val2_749_fu_35976_p2;
wire   [0:0] p_Result_749_fu_35968_p3;
wire   [0:0] p_Result_750_fu_35982_p3;
wire   [0:0] xor_ln895_456_fu_35990_p2;
wire   [0:0] xor_ln896_456_fu_36002_p2;
wire   [0:0] xor_ln302_265_fu_36014_p2;
wire   [0:0] overflow_294_fu_35996_p2;
wire   [0:0] xor_ln302_266_fu_36020_p2;
wire   [0:0] underflow_294_fu_36008_p2;
wire   [0:0] or_ln302_132_fu_36026_p2;
wire   [31:0] select_ln302_265_fu_36032_p3;
wire   [31:0] select_ln350_132_fu_36040_p3;
wire  signed [31:0] lhs_115_fu_35232_p3;
wire  signed [31:0] rhs_133_fu_32331_p3;
wire  signed [32:0] sext_ln813_250_fu_36060_p1;
wire  signed [32:0] sext_ln813_249_fu_36056_p1;
wire   [32:0] ret_V_133_fu_36064_p2;
wire   [31:0] p_Val2_751_fu_36078_p2;
wire   [0:0] p_Result_751_fu_36070_p3;
wire   [0:0] p_Result_752_fu_36084_p3;
wire   [0:0] xor_ln895_457_fu_36092_p2;
wire   [0:0] xor_ln896_457_fu_36104_p2;
wire   [0:0] xor_ln302_267_fu_36116_p2;
wire   [0:0] overflow_295_fu_36098_p2;
wire   [0:0] xor_ln302_268_fu_36122_p2;
wire   [0:0] underflow_295_fu_36110_p2;
wire   [0:0] or_ln302_133_fu_36128_p2;
wire   [31:0] select_ln302_267_fu_36134_p3;
wire   [31:0] select_ln350_133_fu_36142_p3;
wire  signed [31:0] lhs_116_fu_35334_p3;
wire  signed [31:0] rhs_134_fu_32480_p3;
wire  signed [32:0] sext_ln813_252_fu_36162_p1;
wire  signed [32:0] sext_ln813_251_fu_36158_p1;
wire   [32:0] ret_V_134_fu_36166_p2;
wire   [31:0] p_Val2_753_fu_36180_p2;
wire   [0:0] p_Result_753_fu_36172_p3;
wire   [0:0] p_Result_754_fu_36186_p3;
wire   [0:0] xor_ln895_458_fu_36194_p2;
wire   [0:0] xor_ln896_458_fu_36206_p2;
wire   [0:0] xor_ln302_269_fu_36218_p2;
wire   [0:0] overflow_296_fu_36200_p2;
wire   [0:0] xor_ln302_270_fu_36224_p2;
wire   [0:0] underflow_296_fu_36212_p2;
wire   [0:0] or_ln302_134_fu_36230_p2;
wire   [31:0] select_ln302_269_fu_36236_p3;
wire   [31:0] select_ln350_134_fu_36244_p3;
wire  signed [31:0] lhs_117_fu_35436_p3;
wire  signed [31:0] rhs_135_fu_32629_p3;
wire  signed [32:0] sext_ln813_254_fu_36264_p1;
wire  signed [32:0] sext_ln813_253_fu_36260_p1;
wire   [32:0] ret_V_135_fu_36268_p2;
wire   [31:0] p_Val2_755_fu_36282_p2;
wire   [0:0] p_Result_755_fu_36274_p3;
wire   [0:0] p_Result_756_fu_36288_p3;
wire   [0:0] xor_ln895_459_fu_36296_p2;
wire   [0:0] xor_ln896_459_fu_36308_p2;
wire   [0:0] xor_ln302_271_fu_36320_p2;
wire   [0:0] overflow_297_fu_36302_p2;
wire   [0:0] xor_ln302_272_fu_36326_p2;
wire   [0:0] underflow_297_fu_36314_p2;
wire   [0:0] or_ln302_135_fu_36332_p2;
wire   [31:0] select_ln302_271_fu_36338_p3;
wire   [31:0] select_ln350_135_fu_36346_p3;
wire  signed [31:0] lhs_118_fu_35538_p3;
wire  signed [31:0] rhs_136_fu_32778_p3;
wire  signed [32:0] sext_ln813_256_fu_36366_p1;
wire  signed [32:0] sext_ln813_255_fu_36362_p1;
wire   [32:0] ret_V_136_fu_36370_p2;
wire   [31:0] p_Val2_757_fu_36384_p2;
wire   [0:0] p_Result_757_fu_36376_p3;
wire   [0:0] p_Result_758_fu_36390_p3;
wire   [0:0] xor_ln895_460_fu_36398_p2;
wire   [0:0] xor_ln896_460_fu_36410_p2;
wire   [0:0] xor_ln302_273_fu_36422_p2;
wire   [0:0] overflow_298_fu_36404_p2;
wire   [0:0] xor_ln302_274_fu_36428_p2;
wire   [0:0] underflow_298_fu_36416_p2;
wire   [0:0] or_ln302_136_fu_36434_p2;
wire   [31:0] select_ln302_273_fu_36440_p3;
wire   [31:0] select_ln350_136_fu_36448_p3;
wire  signed [31:0] lhs_119_fu_35640_p3;
wire  signed [31:0] rhs_137_fu_32927_p3;
wire  signed [32:0] sext_ln813_258_fu_36468_p1;
wire  signed [32:0] sext_ln813_257_fu_36464_p1;
wire   [32:0] ret_V_137_fu_36472_p2;
wire   [31:0] p_Val2_759_fu_36486_p2;
wire   [0:0] p_Result_759_fu_36478_p3;
wire   [0:0] p_Result_760_fu_36492_p3;
wire   [0:0] xor_ln895_461_fu_36500_p2;
wire   [0:0] xor_ln896_461_fu_36512_p2;
wire   [0:0] xor_ln302_275_fu_36524_p2;
wire   [0:0] overflow_299_fu_36506_p2;
wire   [0:0] xor_ln302_276_fu_36530_p2;
wire   [0:0] underflow_299_fu_36518_p2;
wire   [0:0] or_ln302_137_fu_36536_p2;
wire   [31:0] select_ln302_275_fu_36542_p3;
wire   [31:0] select_ln350_137_fu_36550_p3;
wire  signed [31:0] lhs_120_fu_35742_p3;
wire  signed [31:0] rhs_138_fu_33076_p3;
wire  signed [32:0] sext_ln813_260_fu_36570_p1;
wire  signed [32:0] sext_ln813_259_fu_36566_p1;
wire   [32:0] ret_V_138_fu_36574_p2;
wire   [31:0] p_Val2_761_fu_36588_p2;
wire   [0:0] p_Result_761_fu_36580_p3;
wire   [0:0] p_Result_762_fu_36594_p3;
wire   [0:0] xor_ln895_462_fu_36602_p2;
wire   [0:0] xor_ln896_462_fu_36614_p2;
wire   [0:0] xor_ln302_277_fu_36626_p2;
wire   [0:0] overflow_300_fu_36608_p2;
wire   [0:0] xor_ln302_278_fu_36632_p2;
wire   [0:0] underflow_300_fu_36620_p2;
wire   [0:0] or_ln302_138_fu_36638_p2;
wire   [31:0] select_ln302_277_fu_36644_p3;
wire   [31:0] select_ln350_138_fu_36652_p3;
wire  signed [31:0] lhs_121_fu_35844_p3;
wire  signed [31:0] rhs_139_fu_33225_p3;
wire  signed [32:0] sext_ln813_262_fu_36672_p1;
wire  signed [32:0] sext_ln813_261_fu_36668_p1;
wire   [32:0] ret_V_139_fu_36676_p2;
wire   [31:0] p_Val2_763_fu_36690_p2;
wire   [0:0] p_Result_763_fu_36682_p3;
wire   [0:0] p_Result_764_fu_36696_p3;
wire   [0:0] xor_ln895_463_fu_36704_p2;
wire   [0:0] xor_ln896_463_fu_36716_p2;
wire   [0:0] xor_ln302_279_fu_36728_p2;
wire   [0:0] overflow_301_fu_36710_p2;
wire   [0:0] xor_ln302_280_fu_36734_p2;
wire   [0:0] underflow_301_fu_36722_p2;
wire   [0:0] or_ln302_139_fu_36740_p2;
wire   [31:0] select_ln302_279_fu_36746_p3;
wire   [31:0] select_ln350_139_fu_36754_p3;
wire  signed [31:0] lhs_122_fu_35946_p3;
wire  signed [31:0] rhs_140_fu_33374_p3;
wire  signed [32:0] sext_ln813_264_fu_36774_p1;
wire  signed [32:0] sext_ln813_263_fu_36770_p1;
wire   [32:0] ret_V_140_fu_36778_p2;
wire   [31:0] p_Val2_765_fu_36792_p2;
wire   [0:0] p_Result_765_fu_36784_p3;
wire   [0:0] p_Result_766_fu_36798_p3;
wire   [0:0] xor_ln895_464_fu_36806_p2;
wire   [0:0] xor_ln896_464_fu_36818_p2;
wire   [0:0] xor_ln302_281_fu_36830_p2;
wire   [0:0] overflow_302_fu_36812_p2;
wire   [0:0] xor_ln302_282_fu_36836_p2;
wire   [0:0] underflow_302_fu_36824_p2;
wire   [0:0] or_ln302_140_fu_36842_p2;
wire   [31:0] select_ln302_281_fu_36848_p3;
wire   [31:0] select_ln350_140_fu_36856_p3;
wire  signed [31:0] lhs_123_fu_36048_p3;
wire  signed [31:0] rhs_141_fu_33523_p3;
wire  signed [32:0] sext_ln813_266_fu_36876_p1;
wire  signed [32:0] sext_ln813_265_fu_36872_p1;
wire   [32:0] ret_V_141_fu_36880_p2;
wire   [31:0] p_Val2_767_fu_36894_p2;
wire   [0:0] p_Result_767_fu_36886_p3;
wire   [0:0] p_Result_768_fu_36900_p3;
wire   [0:0] xor_ln895_465_fu_36908_p2;
wire   [0:0] xor_ln896_465_fu_36920_p2;
wire   [0:0] xor_ln302_283_fu_36932_p2;
wire   [0:0] overflow_303_fu_36914_p2;
wire   [0:0] xor_ln302_284_fu_36938_p2;
wire   [0:0] underflow_303_fu_36926_p2;
wire   [0:0] or_ln302_141_fu_36944_p2;
wire   [31:0] select_ln302_283_fu_36950_p3;
wire   [31:0] select_ln350_141_fu_36958_p3;
wire  signed [31:0] lhs_124_fu_36150_p3;
wire  signed [31:0] rhs_142_fu_33541_p3;
wire  signed [32:0] sext_ln813_268_fu_36978_p1;
wire  signed [32:0] sext_ln813_267_fu_36974_p1;
wire   [32:0] ret_V_142_fu_36982_p2;
wire   [31:0] p_Val2_769_fu_36996_p2;
wire   [0:0] p_Result_769_fu_36988_p3;
wire   [0:0] p_Result_770_fu_37002_p3;
wire   [0:0] xor_ln895_466_fu_37010_p2;
wire   [0:0] xor_ln896_466_fu_37022_p2;
wire   [0:0] xor_ln302_285_fu_37034_p2;
wire   [0:0] overflow_304_fu_37016_p2;
wire   [0:0] xor_ln302_286_fu_37040_p2;
wire   [0:0] underflow_304_fu_37028_p2;
wire   [0:0] or_ln302_142_fu_37046_p2;
wire   [31:0] select_ln302_285_fu_37052_p3;
wire   [31:0] select_ln350_142_fu_37060_p3;
wire   [0:0] xor_ln896_368_fu_37076_p2;
wire   [0:0] xor_ln888_284_fu_37086_p2;
wire   [0:0] or_ln888_143_fu_37091_p2;
wire   [0:0] tmp_1020_fu_37101_p3;
wire   [0:0] xor_ln890_141_fu_37109_p2;
wire   [0:0] or_ln890_143_fu_37115_p2;
wire   [0:0] carry_285_fu_37081_p2;
wire   [0:0] deleted_zeros_140_fu_37096_p2;
wire   [0:0] xor_ln895_368_fu_37131_p2;
wire   [0:0] or_ln895_143_fu_37137_p2;
wire   [0:0] xor_ln895_369_fu_37142_p2;
wire   [0:0] deleted_ones_224_fu_37121_p2;
wire   [0:0] xor_ln896_369_fu_37153_p2;
wire   [0:0] and_ln891_143_fu_37126_p2;
wire   [0:0] or_ln896_143_fu_37159_p2;
wire   [0:0] xor_ln896_548_fu_37165_p2;
wire   [0:0] overflow_224_fu_37147_p2;
wire   [0:0] underflow_224_fu_37171_p2;
wire   [0:0] or_ln346_143_fu_37184_p2;
wire   [31:0] select_ln346_225_fu_37176_p3;
wire   [0:0] xor_ln896_370_fu_37200_p2;
wire   [0:0] xor_ln888_286_fu_37210_p2;
wire   [0:0] or_ln888_144_fu_37215_p2;
wire   [0:0] tmp_1026_fu_37225_p3;
wire   [0:0] xor_ln890_142_fu_37233_p2;
wire   [0:0] or_ln890_144_fu_37239_p2;
wire   [0:0] carry_287_fu_37205_p2;
wire   [0:0] deleted_zeros_141_fu_37220_p2;
wire   [0:0] xor_ln895_370_fu_37255_p2;
wire   [0:0] or_ln895_144_fu_37261_p2;
wire   [0:0] xor_ln895_371_fu_37266_p2;
wire   [0:0] deleted_ones_225_fu_37245_p2;
wire   [0:0] xor_ln896_371_fu_37277_p2;
wire   [0:0] and_ln891_144_fu_37250_p2;
wire   [0:0] or_ln896_144_fu_37283_p2;
wire   [0:0] xor_ln896_549_fu_37289_p2;
wire   [0:0] overflow_225_fu_37271_p2;
wire   [0:0] underflow_225_fu_37295_p2;
wire   [0:0] or_ln346_144_fu_37308_p2;
wire   [31:0] select_ln346_226_fu_37300_p3;
wire  signed [31:0] sext_ln856_137_fu_37197_p1;
wire   [0:0] xor_ln896_372_fu_37325_p2;
wire   [0:0] xor_ln888_288_fu_37335_p2;
wire   [0:0] or_ln888_145_fu_37340_p2;
wire   [0:0] tmp_1032_fu_37350_p3;
wire   [0:0] xor_ln890_143_fu_37358_p2;
wire   [0:0] or_ln890_145_fu_37364_p2;
wire   [0:0] carry_289_fu_37330_p2;
wire   [0:0] deleted_zeros_142_fu_37345_p2;
wire   [0:0] xor_ln895_372_fu_37380_p2;
wire   [0:0] or_ln895_145_fu_37386_p2;
wire   [0:0] xor_ln895_373_fu_37391_p2;
wire   [0:0] deleted_ones_226_fu_37370_p2;
wire   [0:0] xor_ln896_373_fu_37402_p2;
wire   [0:0] and_ln891_145_fu_37375_p2;
wire   [0:0] or_ln896_145_fu_37408_p2;
wire   [0:0] xor_ln896_550_fu_37414_p2;
wire   [0:0] overflow_226_fu_37396_p2;
wire   [0:0] underflow_226_fu_37420_p2;
wire   [0:0] or_ln346_145_fu_37433_p2;
wire   [31:0] select_ln346_227_fu_37425_p3;
wire  signed [31:0] sext_ln856_138_fu_37322_p1;
wire   [0:0] xor_ln896_374_fu_37450_p2;
wire   [0:0] xor_ln888_290_fu_37460_p2;
wire   [0:0] or_ln888_146_fu_37465_p2;
wire   [0:0] tmp_1038_fu_37475_p3;
wire   [0:0] xor_ln890_144_fu_37483_p2;
wire   [0:0] or_ln890_146_fu_37489_p2;
wire   [0:0] carry_291_fu_37455_p2;
wire   [0:0] deleted_zeros_143_fu_37470_p2;
wire   [0:0] xor_ln895_374_fu_37505_p2;
wire   [0:0] or_ln895_146_fu_37511_p2;
wire   [0:0] xor_ln895_375_fu_37516_p2;
wire   [0:0] deleted_ones_227_fu_37495_p2;
wire   [0:0] xor_ln896_375_fu_37527_p2;
wire   [0:0] and_ln891_146_fu_37500_p2;
wire   [0:0] or_ln896_146_fu_37533_p2;
wire   [0:0] xor_ln896_551_fu_37539_p2;
wire   [0:0] overflow_227_fu_37521_p2;
wire   [0:0] underflow_227_fu_37545_p2;
wire   [0:0] or_ln346_146_fu_37558_p2;
wire   [31:0] select_ln346_228_fu_37550_p3;
wire  signed [31:0] sext_ln856_139_fu_37447_p1;
wire   [0:0] xor_ln896_376_fu_37575_p2;
wire   [0:0] xor_ln888_292_fu_37585_p2;
wire   [0:0] or_ln888_147_fu_37590_p2;
wire   [0:0] tmp_1044_fu_37600_p3;
wire   [0:0] xor_ln890_145_fu_37608_p2;
wire   [0:0] or_ln890_147_fu_37614_p2;
wire   [0:0] carry_293_fu_37580_p2;
wire   [0:0] deleted_zeros_144_fu_37595_p2;
wire   [0:0] xor_ln895_376_fu_37630_p2;
wire   [0:0] or_ln895_147_fu_37636_p2;
wire   [0:0] xor_ln895_377_fu_37641_p2;
wire   [0:0] deleted_ones_228_fu_37620_p2;
wire   [0:0] xor_ln896_377_fu_37652_p2;
wire   [0:0] and_ln891_147_fu_37625_p2;
wire   [0:0] or_ln896_147_fu_37658_p2;
wire   [0:0] xor_ln896_552_fu_37664_p2;
wire   [0:0] overflow_228_fu_37646_p2;
wire   [0:0] underflow_228_fu_37670_p2;
wire   [0:0] or_ln346_147_fu_37683_p2;
wire   [31:0] select_ln346_229_fu_37675_p3;
wire  signed [31:0] sext_ln856_140_fu_37572_p1;
wire   [0:0] xor_ln896_378_fu_37700_p2;
wire   [0:0] xor_ln888_294_fu_37710_p2;
wire   [0:0] or_ln888_148_fu_37715_p2;
wire   [0:0] tmp_1050_fu_37725_p3;
wire   [0:0] xor_ln890_146_fu_37733_p2;
wire   [0:0] or_ln890_148_fu_37739_p2;
wire   [0:0] carry_295_fu_37705_p2;
wire   [0:0] deleted_zeros_145_fu_37720_p2;
wire   [0:0] xor_ln895_378_fu_37755_p2;
wire   [0:0] or_ln895_148_fu_37761_p2;
wire   [0:0] xor_ln895_379_fu_37766_p2;
wire   [0:0] deleted_ones_229_fu_37745_p2;
wire   [0:0] xor_ln896_379_fu_37777_p2;
wire   [0:0] and_ln891_148_fu_37750_p2;
wire   [0:0] or_ln896_148_fu_37783_p2;
wire   [0:0] xor_ln896_553_fu_37789_p2;
wire   [0:0] overflow_229_fu_37771_p2;
wire   [0:0] underflow_229_fu_37795_p2;
wire   [0:0] or_ln346_148_fu_37808_p2;
wire   [31:0] select_ln346_230_fu_37800_p3;
wire  signed [31:0] sext_ln856_141_fu_37697_p1;
wire   [0:0] xor_ln896_380_fu_37825_p2;
wire   [0:0] xor_ln888_296_fu_37835_p2;
wire   [0:0] or_ln888_149_fu_37840_p2;
wire   [0:0] tmp_1056_fu_37850_p3;
wire   [0:0] xor_ln890_147_fu_37858_p2;
wire   [0:0] or_ln890_149_fu_37864_p2;
wire   [0:0] carry_297_fu_37830_p2;
wire   [0:0] deleted_zeros_146_fu_37845_p2;
wire   [0:0] xor_ln895_380_fu_37880_p2;
wire   [0:0] or_ln895_149_fu_37886_p2;
wire   [0:0] xor_ln895_381_fu_37891_p2;
wire   [0:0] deleted_ones_230_fu_37870_p2;
wire   [0:0] xor_ln896_381_fu_37902_p2;
wire   [0:0] and_ln891_149_fu_37875_p2;
wire   [0:0] or_ln896_149_fu_37908_p2;
wire   [0:0] xor_ln896_554_fu_37914_p2;
wire   [0:0] overflow_230_fu_37896_p2;
wire   [0:0] underflow_230_fu_37920_p2;
wire   [0:0] or_ln346_149_fu_37933_p2;
wire   [31:0] select_ln346_231_fu_37925_p3;
wire  signed [31:0] sext_ln856_142_fu_37822_p1;
wire   [0:0] xor_ln896_382_fu_37950_p2;
wire   [0:0] xor_ln888_298_fu_37960_p2;
wire   [0:0] or_ln888_150_fu_37965_p2;
wire   [0:0] tmp_1062_fu_37975_p3;
wire   [0:0] xor_ln890_148_fu_37983_p2;
wire   [0:0] or_ln890_150_fu_37989_p2;
wire   [0:0] carry_299_fu_37955_p2;
wire   [0:0] deleted_zeros_147_fu_37970_p2;
wire   [0:0] xor_ln895_382_fu_38005_p2;
wire   [0:0] or_ln895_150_fu_38011_p2;
wire   [0:0] xor_ln895_383_fu_38016_p2;
wire   [0:0] deleted_ones_231_fu_37995_p2;
wire   [0:0] xor_ln896_383_fu_38027_p2;
wire   [0:0] and_ln891_150_fu_38000_p2;
wire   [0:0] or_ln896_150_fu_38033_p2;
wire   [0:0] xor_ln896_555_fu_38039_p2;
wire   [0:0] overflow_231_fu_38021_p2;
wire   [0:0] underflow_231_fu_38045_p2;
wire   [0:0] or_ln346_150_fu_38058_p2;
wire   [31:0] select_ln346_232_fu_38050_p3;
wire  signed [31:0] sext_ln856_143_fu_37947_p1;
wire   [0:0] xor_ln896_384_fu_38075_p2;
wire   [0:0] xor_ln888_300_fu_38085_p2;
wire   [0:0] or_ln888_151_fu_38090_p2;
wire   [0:0] tmp_1068_fu_38100_p3;
wire   [0:0] xor_ln890_149_fu_38108_p2;
wire   [0:0] or_ln890_151_fu_38114_p2;
wire   [0:0] carry_301_fu_38080_p2;
wire   [0:0] deleted_zeros_148_fu_38095_p2;
wire   [0:0] xor_ln895_384_fu_38130_p2;
wire   [0:0] or_ln895_151_fu_38136_p2;
wire   [0:0] xor_ln895_385_fu_38141_p2;
wire   [0:0] deleted_ones_232_fu_38120_p2;
wire   [0:0] xor_ln896_385_fu_38152_p2;
wire   [0:0] and_ln891_151_fu_38125_p2;
wire   [0:0] or_ln896_151_fu_38158_p2;
wire   [0:0] xor_ln896_556_fu_38164_p2;
wire   [0:0] overflow_232_fu_38146_p2;
wire   [0:0] underflow_232_fu_38170_p2;
wire   [0:0] or_ln346_151_fu_38183_p2;
wire   [31:0] select_ln346_233_fu_38175_p3;
wire  signed [31:0] sext_ln856_144_fu_38072_p1;
wire   [31:0] zext_ln377_152_fu_38200_p1;
wire  signed [31:0] sext_ln818_3_fu_38197_p1;
wire   [31:0] p_Val2_619_fu_38203_p2;
wire   [0:0] p_Result_620_fu_38209_p3;
wire   [0:0] xor_ln896_386_fu_38217_p2;
wire   [0:0] xor_ln888_302_fu_38228_p2;
wire   [0:0] or_ln888_152_fu_38233_p2;
wire   [0:0] tmp_1074_fu_38244_p3;
wire   [0:0] xor_ln890_150_fu_38252_p2;
wire   [0:0] or_ln890_152_fu_38258_p2;
wire   [0:0] carry_303_fu_38223_p2;
wire   [0:0] deleted_zeros_149_fu_38239_p2;
wire   [0:0] xor_ln895_386_fu_38274_p2;
wire   [0:0] or_ln895_152_fu_38280_p2;
wire   [0:0] xor_ln895_387_fu_38286_p2;
wire   [0:0] deleted_ones_233_fu_38264_p2;
wire   [0:0] xor_ln896_387_fu_38297_p2;
wire   [0:0] and_ln891_152_fu_38269_p2;
wire   [0:0] or_ln896_152_fu_38303_p2;
wire   [0:0] xor_ln896_557_fu_38309_p2;
wire   [0:0] overflow_233_fu_38291_p2;
wire   [0:0] underflow_233_fu_38315_p2;
wire   [0:0] or_ln346_152_fu_38328_p2;
wire   [31:0] select_ln346_234_fu_38320_p3;
wire   [18:0] zext_ln377_153_fu_38345_p1;
wire  signed [18:0] sext_ln823_145_fu_38342_p1;
wire  signed [18:0] p_Val2_622_fu_38348_p2;
wire   [0:0] p_Result_623_fu_38358_p3;
wire   [0:0] xor_ln896_388_fu_38366_p2;
wire   [0:0] xor_ln888_304_fu_38377_p2;
wire   [0:0] or_ln888_153_fu_38382_p2;
wire   [0:0] tmp_1080_fu_38393_p3;
wire   [0:0] xor_ln890_151_fu_38401_p2;
wire   [0:0] or_ln890_153_fu_38407_p2;
wire   [0:0] carry_305_fu_38372_p2;
wire   [0:0] deleted_zeros_150_fu_38388_p2;
wire   [0:0] xor_ln895_388_fu_38423_p2;
wire   [0:0] or_ln895_153_fu_38429_p2;
wire   [0:0] xor_ln895_389_fu_38435_p2;
wire   [0:0] deleted_ones_234_fu_38413_p2;
wire   [0:0] xor_ln896_389_fu_38446_p2;
wire   [0:0] and_ln891_153_fu_38418_p2;
wire   [0:0] or_ln896_153_fu_38452_p2;
wire   [0:0] xor_ln896_558_fu_38458_p2;
wire   [0:0] overflow_234_fu_38440_p2;
wire   [0:0] underflow_234_fu_38464_p2;
wire   [0:0] or_ln346_153_fu_38477_p2;
wire   [31:0] select_ln346_235_fu_38469_p3;
wire  signed [31:0] sext_ln856_145_fu_38354_p1;
wire   [20:0] zext_ln377_154_fu_38494_p1;
wire  signed [20:0] sext_ln823_146_fu_38491_p1;
wire  signed [20:0] p_Val2_625_fu_38497_p2;
wire   [0:0] p_Result_626_fu_38507_p3;
wire   [0:0] xor_ln896_390_fu_38515_p2;
wire   [0:0] xor_ln888_306_fu_38526_p2;
wire   [0:0] or_ln888_154_fu_38531_p2;
wire   [0:0] tmp_1086_fu_38542_p3;
wire   [0:0] xor_ln890_152_fu_38550_p2;
wire   [0:0] or_ln890_154_fu_38556_p2;
wire   [0:0] carry_307_fu_38521_p2;
wire   [0:0] deleted_zeros_151_fu_38537_p2;
wire   [0:0] xor_ln895_390_fu_38572_p2;
wire   [0:0] or_ln895_154_fu_38578_p2;
wire   [0:0] xor_ln895_391_fu_38584_p2;
wire   [0:0] deleted_ones_235_fu_38562_p2;
wire   [0:0] xor_ln896_391_fu_38595_p2;
wire   [0:0] and_ln891_154_fu_38567_p2;
wire   [0:0] or_ln896_154_fu_38601_p2;
wire   [0:0] xor_ln896_559_fu_38607_p2;
wire   [0:0] overflow_235_fu_38589_p2;
wire   [0:0] underflow_235_fu_38613_p2;
wire   [0:0] or_ln346_154_fu_38626_p2;
wire   [31:0] select_ln346_236_fu_38618_p3;
wire  signed [31:0] sext_ln856_146_fu_38503_p1;
wire   [26:0] zext_ln377_155_fu_38643_p1;
wire  signed [26:0] sext_ln823_147_fu_38640_p1;
wire  signed [26:0] p_Val2_628_fu_38646_p2;
wire   [0:0] p_Result_629_fu_38656_p3;
wire   [0:0] xor_ln896_392_fu_38664_p2;
wire   [0:0] xor_ln888_308_fu_38675_p2;
wire   [0:0] or_ln888_155_fu_38680_p2;
wire   [0:0] tmp_1092_fu_38691_p3;
wire   [0:0] xor_ln890_153_fu_38699_p2;
wire   [0:0] or_ln890_155_fu_38705_p2;
wire   [0:0] carry_309_fu_38670_p2;
wire   [0:0] deleted_zeros_152_fu_38686_p2;
wire   [0:0] xor_ln895_392_fu_38721_p2;
wire   [0:0] or_ln895_155_fu_38727_p2;
wire   [0:0] xor_ln895_393_fu_38733_p2;
wire   [0:0] deleted_ones_236_fu_38711_p2;
wire   [0:0] xor_ln896_393_fu_38744_p2;
wire   [0:0] and_ln891_155_fu_38716_p2;
wire   [0:0] or_ln896_155_fu_38750_p2;
wire   [0:0] xor_ln896_560_fu_38756_p2;
wire   [0:0] overflow_236_fu_38738_p2;
wire   [0:0] underflow_236_fu_38762_p2;
wire   [0:0] or_ln346_155_fu_38775_p2;
wire   [31:0] select_ln346_237_fu_38767_p3;
wire  signed [31:0] sext_ln856_147_fu_38652_p1;
wire   [26:0] zext_ln377_156_fu_38792_p1;
wire  signed [26:0] sext_ln823_148_fu_38789_p1;
wire  signed [26:0] p_Val2_631_fu_38795_p2;
wire   [0:0] p_Result_632_fu_38805_p3;
wire   [0:0] xor_ln896_394_fu_38813_p2;
wire   [0:0] xor_ln888_310_fu_38824_p2;
wire   [0:0] or_ln888_156_fu_38829_p2;
wire   [0:0] tmp_1098_fu_38840_p3;
wire   [0:0] xor_ln890_154_fu_38848_p2;
wire   [0:0] or_ln890_156_fu_38854_p2;
wire   [0:0] carry_311_fu_38819_p2;
wire   [0:0] deleted_zeros_153_fu_38835_p2;
wire   [0:0] xor_ln895_394_fu_38870_p2;
wire   [0:0] or_ln895_156_fu_38876_p2;
wire   [0:0] xor_ln895_395_fu_38882_p2;
wire   [0:0] deleted_ones_237_fu_38860_p2;
wire   [0:0] xor_ln896_395_fu_38893_p2;
wire   [0:0] and_ln891_156_fu_38865_p2;
wire   [0:0] or_ln896_156_fu_38899_p2;
wire   [0:0] xor_ln896_561_fu_38905_p2;
wire   [0:0] overflow_237_fu_38887_p2;
wire   [0:0] underflow_237_fu_38911_p2;
wire   [0:0] or_ln346_156_fu_38924_p2;
wire   [31:0] select_ln346_238_fu_38916_p3;
wire  signed [31:0] sext_ln856_148_fu_38801_p1;
wire   [18:0] zext_ln377_157_fu_38941_p1;
wire  signed [18:0] sext_ln823_149_fu_38938_p1;
wire  signed [18:0] p_Val2_634_fu_38944_p2;
wire   [0:0] p_Result_635_fu_38954_p3;
wire   [0:0] xor_ln896_396_fu_38962_p2;
wire   [0:0] xor_ln888_312_fu_38973_p2;
wire   [0:0] or_ln888_157_fu_38978_p2;
wire   [0:0] tmp_1104_fu_38989_p3;
wire   [0:0] xor_ln890_155_fu_38997_p2;
wire   [0:0] or_ln890_157_fu_39003_p2;
wire   [0:0] carry_313_fu_38968_p2;
wire   [0:0] deleted_zeros_154_fu_38984_p2;
wire   [0:0] xor_ln895_396_fu_39019_p2;
wire   [0:0] or_ln895_157_fu_39025_p2;
wire   [0:0] xor_ln895_397_fu_39031_p2;
wire   [0:0] deleted_ones_238_fu_39009_p2;
wire   [0:0] xor_ln896_397_fu_39042_p2;
wire   [0:0] and_ln891_157_fu_39014_p2;
wire   [0:0] or_ln896_157_fu_39048_p2;
wire   [0:0] xor_ln896_562_fu_39054_p2;
wire   [0:0] overflow_238_fu_39036_p2;
wire   [0:0] underflow_238_fu_39060_p2;
wire   [0:0] or_ln346_157_fu_39073_p2;
wire   [31:0] select_ln346_239_fu_39065_p3;
wire  signed [31:0] sext_ln856_149_fu_38950_p1;
wire   [20:0] zext_ln377_158_fu_39090_p1;
wire  signed [20:0] sext_ln823_150_fu_39087_p1;
wire  signed [20:0] p_Val2_637_fu_39093_p2;
wire   [0:0] p_Result_638_fu_39103_p3;
wire   [0:0] xor_ln896_398_fu_39111_p2;
wire   [0:0] xor_ln888_314_fu_39122_p2;
wire   [0:0] or_ln888_158_fu_39127_p2;
wire   [0:0] tmp_1110_fu_39138_p3;
wire   [0:0] xor_ln890_156_fu_39146_p2;
wire   [0:0] or_ln890_158_fu_39152_p2;
wire   [0:0] carry_315_fu_39117_p2;
wire   [0:0] deleted_zeros_155_fu_39133_p2;
wire   [0:0] xor_ln895_398_fu_39168_p2;
wire   [0:0] or_ln895_158_fu_39174_p2;
wire   [0:0] xor_ln895_399_fu_39180_p2;
wire   [0:0] deleted_ones_239_fu_39158_p2;
wire   [0:0] xor_ln896_399_fu_39191_p2;
wire   [0:0] and_ln891_158_fu_39163_p2;
wire   [0:0] or_ln896_158_fu_39197_p2;
wire   [0:0] xor_ln896_563_fu_39203_p2;
wire   [0:0] overflow_239_fu_39185_p2;
wire   [0:0] underflow_239_fu_39209_p2;
wire   [0:0] or_ln346_158_fu_39222_p2;
wire   [31:0] select_ln346_240_fu_39214_p3;
wire  signed [31:0] sext_ln856_150_fu_39099_p1;
wire   [31:0] select_ln346_241_fu_39239_p3;
wire  signed [31:0] sext_ln856_151_fu_39236_p1;
wire   [26:0] zext_ln377_160_fu_39256_p1;
wire  signed [26:0] sext_ln823_152_fu_39253_p1;
wire  signed [26:0] p_Val2_643_fu_39259_p2;
wire   [0:0] p_Result_644_fu_39269_p3;
wire   [0:0] xor_ln896_402_fu_39277_p2;
wire   [0:0] xor_ln888_318_fu_39288_p2;
wire   [0:0] or_ln888_160_fu_39293_p2;
wire   [0:0] tmp_1122_fu_39304_p3;
wire   [0:0] xor_ln890_158_fu_39312_p2;
wire   [0:0] or_ln890_160_fu_39318_p2;
wire   [0:0] carry_319_fu_39283_p2;
wire   [0:0] deleted_zeros_157_fu_39299_p2;
wire   [0:0] xor_ln895_402_fu_39334_p2;
wire   [0:0] or_ln895_160_fu_39340_p2;
wire   [0:0] xor_ln895_403_fu_39346_p2;
wire   [0:0] deleted_ones_241_fu_39324_p2;
wire   [0:0] xor_ln896_403_fu_39357_p2;
wire   [0:0] and_ln891_160_fu_39329_p2;
wire   [0:0] or_ln896_160_fu_39363_p2;
wire   [0:0] xor_ln896_565_fu_39369_p2;
wire   [0:0] overflow_241_fu_39351_p2;
wire   [0:0] underflow_241_fu_39375_p2;
wire   [0:0] or_ln346_160_fu_39388_p2;
wire   [31:0] select_ln346_242_fu_39380_p3;
wire  signed [31:0] sext_ln856_152_fu_39265_p1;
wire  signed [31:0] rhs_143_fu_37190_p3;
wire  signed [32:0] sext_ln813_270_fu_39405_p1;
wire  signed [32:0] sext_ln813_269_fu_39402_p1;
wire   [32:0] ret_V_143_fu_39409_p2;
wire   [31:0] p_Val2_771_fu_39423_p2;
wire   [0:0] p_Result_771_fu_39415_p3;
wire   [0:0] p_Result_772_fu_39428_p3;
wire   [0:0] xor_ln895_467_fu_39436_p2;
wire   [0:0] xor_ln896_467_fu_39448_p2;
wire   [0:0] xor_ln302_287_fu_39460_p2;
wire   [0:0] overflow_305_fu_39442_p2;
wire   [0:0] xor_ln302_288_fu_39466_p2;
wire   [0:0] underflow_305_fu_39454_p2;
wire   [0:0] or_ln302_143_fu_39472_p2;
wire   [31:0] select_ln302_287_fu_39478_p3;
wire   [31:0] select_ln350_143_fu_39486_p3;
wire  signed [31:0] rhs_144_fu_37314_p3;
wire  signed [32:0] sext_ln813_272_fu_39505_p1;
wire  signed [32:0] sext_ln813_271_fu_39502_p1;
wire   [32:0] ret_V_144_fu_39509_p2;
wire   [31:0] p_Val2_773_fu_39523_p2;
wire   [0:0] p_Result_773_fu_39515_p3;
wire   [0:0] p_Result_774_fu_39528_p3;
wire   [0:0] xor_ln895_468_fu_39536_p2;
wire   [0:0] xor_ln896_468_fu_39548_p2;
wire   [0:0] xor_ln302_289_fu_39560_p2;
wire   [0:0] overflow_306_fu_39542_p2;
wire   [0:0] xor_ln302_290_fu_39566_p2;
wire   [0:0] underflow_306_fu_39554_p2;
wire   [0:0] or_ln302_144_fu_39572_p2;
wire   [31:0] select_ln302_289_fu_39578_p3;
wire   [31:0] select_ln350_144_fu_39586_p3;
wire  signed [31:0] rhs_145_fu_37439_p3;
wire  signed [32:0] sext_ln813_274_fu_39605_p1;
wire  signed [32:0] sext_ln813_273_fu_39602_p1;
wire   [32:0] ret_V_145_fu_39609_p2;
wire   [31:0] p_Val2_775_fu_39623_p2;
wire   [0:0] p_Result_775_fu_39615_p3;
wire   [0:0] p_Result_776_fu_39628_p3;
wire   [0:0] xor_ln895_469_fu_39636_p2;
wire   [0:0] xor_ln896_469_fu_39648_p2;
wire   [0:0] xor_ln302_291_fu_39660_p2;
wire   [0:0] overflow_307_fu_39642_p2;
wire   [0:0] xor_ln302_292_fu_39666_p2;
wire   [0:0] underflow_307_fu_39654_p2;
wire   [0:0] or_ln302_145_fu_39672_p2;
wire   [31:0] select_ln302_291_fu_39678_p3;
wire   [31:0] select_ln350_145_fu_39686_p3;
wire  signed [31:0] rhs_146_fu_37564_p3;
wire  signed [32:0] sext_ln813_276_fu_39705_p1;
wire  signed [32:0] sext_ln813_275_fu_39702_p1;
wire   [32:0] ret_V_146_fu_39709_p2;
wire   [31:0] p_Val2_777_fu_39723_p2;
wire   [0:0] p_Result_777_fu_39715_p3;
wire   [0:0] p_Result_778_fu_39728_p3;
wire   [0:0] xor_ln895_470_fu_39736_p2;
wire   [0:0] xor_ln896_470_fu_39748_p2;
wire   [0:0] xor_ln302_293_fu_39760_p2;
wire   [0:0] overflow_308_fu_39742_p2;
wire   [0:0] xor_ln302_294_fu_39766_p2;
wire   [0:0] underflow_308_fu_39754_p2;
wire   [0:0] or_ln302_146_fu_39772_p2;
wire   [31:0] select_ln302_293_fu_39778_p3;
wire   [31:0] select_ln350_146_fu_39786_p3;
wire  signed [31:0] rhs_147_fu_37689_p3;
wire  signed [32:0] sext_ln813_278_fu_39805_p1;
wire  signed [32:0] sext_ln813_277_fu_39802_p1;
wire   [32:0] ret_V_147_fu_39809_p2;
wire   [31:0] p_Val2_779_fu_39823_p2;
wire   [0:0] p_Result_779_fu_39815_p3;
wire   [0:0] p_Result_780_fu_39828_p3;
wire   [0:0] xor_ln895_471_fu_39836_p2;
wire   [0:0] xor_ln896_471_fu_39848_p2;
wire   [0:0] xor_ln302_295_fu_39860_p2;
wire   [0:0] overflow_309_fu_39842_p2;
wire   [0:0] xor_ln302_296_fu_39866_p2;
wire   [0:0] underflow_309_fu_39854_p2;
wire   [0:0] or_ln302_147_fu_39872_p2;
wire   [31:0] select_ln302_295_fu_39878_p3;
wire   [31:0] select_ln350_147_fu_39886_p3;
wire  signed [31:0] rhs_148_fu_37814_p3;
wire  signed [32:0] sext_ln813_280_fu_39905_p1;
wire  signed [32:0] sext_ln813_279_fu_39902_p1;
wire   [32:0] ret_V_148_fu_39909_p2;
wire   [31:0] p_Val2_781_fu_39923_p2;
wire   [0:0] p_Result_781_fu_39915_p3;
wire   [0:0] p_Result_782_fu_39928_p3;
wire   [0:0] xor_ln895_472_fu_39936_p2;
wire   [0:0] xor_ln896_472_fu_39948_p2;
wire   [0:0] xor_ln302_297_fu_39960_p2;
wire   [0:0] overflow_310_fu_39942_p2;
wire   [0:0] xor_ln302_298_fu_39966_p2;
wire   [0:0] underflow_310_fu_39954_p2;
wire   [0:0] or_ln302_148_fu_39972_p2;
wire   [31:0] select_ln302_297_fu_39978_p3;
wire   [31:0] select_ln350_148_fu_39986_p3;
wire  signed [31:0] rhs_149_fu_37939_p3;
wire  signed [32:0] sext_ln813_282_fu_40005_p1;
wire  signed [32:0] sext_ln813_281_fu_40002_p1;
wire   [32:0] ret_V_149_fu_40009_p2;
wire   [31:0] p_Val2_783_fu_40023_p2;
wire   [0:0] p_Result_783_fu_40015_p3;
wire   [0:0] p_Result_784_fu_40028_p3;
wire   [0:0] xor_ln895_473_fu_40036_p2;
wire   [0:0] xor_ln896_473_fu_40048_p2;
wire   [0:0] xor_ln302_299_fu_40060_p2;
wire   [0:0] overflow_311_fu_40042_p2;
wire   [0:0] xor_ln302_300_fu_40066_p2;
wire   [0:0] underflow_311_fu_40054_p2;
wire   [0:0] or_ln302_149_fu_40072_p2;
wire   [31:0] select_ln302_299_fu_40078_p3;
wire   [31:0] select_ln350_149_fu_40086_p3;
wire  signed [31:0] rhs_150_fu_38064_p3;
wire  signed [32:0] sext_ln813_284_fu_40105_p1;
wire  signed [32:0] sext_ln813_283_fu_40102_p1;
wire   [32:0] ret_V_150_fu_40109_p2;
wire   [31:0] p_Val2_785_fu_40123_p2;
wire   [0:0] p_Result_785_fu_40115_p3;
wire   [0:0] p_Result_786_fu_40128_p3;
wire   [0:0] xor_ln895_474_fu_40136_p2;
wire   [0:0] xor_ln896_474_fu_40148_p2;
wire   [0:0] xor_ln302_301_fu_40160_p2;
wire   [0:0] overflow_312_fu_40142_p2;
wire   [0:0] xor_ln302_302_fu_40166_p2;
wire   [0:0] underflow_312_fu_40154_p2;
wire   [0:0] or_ln302_150_fu_40172_p2;
wire   [31:0] select_ln302_301_fu_40178_p3;
wire   [31:0] select_ln350_150_fu_40186_p3;
wire  signed [31:0] rhs_151_fu_38189_p3;
wire  signed [32:0] sext_ln813_286_fu_40205_p1;
wire  signed [32:0] sext_ln813_285_fu_40202_p1;
wire   [32:0] ret_V_151_fu_40209_p2;
wire   [31:0] p_Val2_787_fu_40223_p2;
wire   [0:0] p_Result_787_fu_40215_p3;
wire   [0:0] p_Result_788_fu_40228_p3;
wire   [0:0] xor_ln895_475_fu_40236_p2;
wire   [0:0] xor_ln896_475_fu_40248_p2;
wire   [0:0] xor_ln302_303_fu_40260_p2;
wire   [0:0] overflow_313_fu_40242_p2;
wire   [0:0] xor_ln302_304_fu_40266_p2;
wire   [0:0] underflow_313_fu_40254_p2;
wire   [0:0] or_ln302_151_fu_40272_p2;
wire   [31:0] select_ln302_303_fu_40278_p3;
wire   [31:0] select_ln350_151_fu_40286_p3;
wire  signed [31:0] lhs_134_fu_39494_p3;
wire  signed [31:0] rhs_152_fu_38334_p3;
wire  signed [32:0] sext_ln813_288_fu_40306_p1;
wire  signed [32:0] sext_ln813_287_fu_40302_p1;
wire   [32:0] ret_V_152_fu_40310_p2;
wire   [31:0] p_Val2_789_fu_40324_p2;
wire   [0:0] p_Result_789_fu_40316_p3;
wire   [0:0] p_Result_790_fu_40330_p3;
wire   [0:0] xor_ln895_476_fu_40338_p2;
wire   [0:0] xor_ln896_476_fu_40350_p2;
wire   [0:0] xor_ln302_305_fu_40362_p2;
wire   [0:0] overflow_314_fu_40344_p2;
wire   [0:0] xor_ln302_306_fu_40368_p2;
wire   [0:0] underflow_314_fu_40356_p2;
wire   [0:0] or_ln302_152_fu_40374_p2;
wire   [31:0] select_ln302_305_fu_40380_p3;
wire   [31:0] select_ln350_152_fu_40388_p3;
wire  signed [31:0] lhs_135_fu_39594_p3;
wire  signed [31:0] rhs_153_fu_38483_p3;
wire  signed [32:0] sext_ln813_290_fu_40408_p1;
wire  signed [32:0] sext_ln813_289_fu_40404_p1;
wire   [32:0] ret_V_153_fu_40412_p2;
wire   [31:0] p_Val2_791_fu_40426_p2;
wire   [0:0] p_Result_791_fu_40418_p3;
wire   [0:0] p_Result_792_fu_40432_p3;
wire   [0:0] xor_ln895_477_fu_40440_p2;
wire   [0:0] xor_ln896_477_fu_40452_p2;
wire   [0:0] xor_ln302_307_fu_40464_p2;
wire   [0:0] overflow_315_fu_40446_p2;
wire   [0:0] xor_ln302_308_fu_40470_p2;
wire   [0:0] underflow_315_fu_40458_p2;
wire   [0:0] or_ln302_153_fu_40476_p2;
wire   [31:0] select_ln302_307_fu_40482_p3;
wire   [31:0] select_ln350_153_fu_40490_p3;
wire  signed [31:0] lhs_136_fu_39694_p3;
wire  signed [31:0] rhs_154_fu_38632_p3;
wire  signed [32:0] sext_ln813_292_fu_40510_p1;
wire  signed [32:0] sext_ln813_291_fu_40506_p1;
wire   [32:0] ret_V_154_fu_40514_p2;
wire   [31:0] p_Val2_793_fu_40528_p2;
wire   [0:0] p_Result_793_fu_40520_p3;
wire   [0:0] p_Result_794_fu_40534_p3;
wire   [0:0] xor_ln895_478_fu_40542_p2;
wire   [0:0] xor_ln896_478_fu_40554_p2;
wire   [0:0] xor_ln302_309_fu_40566_p2;
wire   [0:0] overflow_316_fu_40548_p2;
wire   [0:0] xor_ln302_310_fu_40572_p2;
wire   [0:0] underflow_316_fu_40560_p2;
wire   [0:0] or_ln302_154_fu_40578_p2;
wire   [31:0] select_ln302_309_fu_40584_p3;
wire   [31:0] select_ln350_154_fu_40592_p3;
wire  signed [31:0] lhs_137_fu_39794_p3;
wire  signed [31:0] rhs_155_fu_38781_p3;
wire  signed [32:0] sext_ln813_294_fu_40612_p1;
wire  signed [32:0] sext_ln813_293_fu_40608_p1;
wire   [32:0] ret_V_155_fu_40616_p2;
wire   [31:0] p_Val2_795_fu_40630_p2;
wire   [0:0] p_Result_795_fu_40622_p3;
wire   [0:0] p_Result_796_fu_40636_p3;
wire   [0:0] xor_ln895_479_fu_40644_p2;
wire   [0:0] xor_ln896_479_fu_40656_p2;
wire   [0:0] xor_ln302_311_fu_40668_p2;
wire   [0:0] overflow_317_fu_40650_p2;
wire   [0:0] xor_ln302_312_fu_40674_p2;
wire   [0:0] underflow_317_fu_40662_p2;
wire   [0:0] or_ln302_155_fu_40680_p2;
wire   [31:0] select_ln302_311_fu_40686_p3;
wire   [31:0] select_ln350_155_fu_40694_p3;
wire  signed [31:0] lhs_138_fu_39894_p3;
wire  signed [31:0] rhs_156_fu_38930_p3;
wire  signed [32:0] sext_ln813_296_fu_40714_p1;
wire  signed [32:0] sext_ln813_295_fu_40710_p1;
wire   [32:0] ret_V_156_fu_40718_p2;
wire   [31:0] p_Val2_797_fu_40732_p2;
wire   [0:0] p_Result_797_fu_40724_p3;
wire   [0:0] p_Result_798_fu_40738_p3;
wire   [0:0] xor_ln895_480_fu_40746_p2;
wire   [0:0] xor_ln896_480_fu_40758_p2;
wire   [0:0] xor_ln302_313_fu_40770_p2;
wire   [0:0] overflow_318_fu_40752_p2;
wire   [0:0] xor_ln302_314_fu_40776_p2;
wire   [0:0] underflow_318_fu_40764_p2;
wire   [0:0] or_ln302_156_fu_40782_p2;
wire   [31:0] select_ln302_313_fu_40788_p3;
wire   [31:0] select_ln350_156_fu_40796_p3;
wire  signed [31:0] lhs_139_fu_39994_p3;
wire  signed [31:0] rhs_157_fu_39079_p3;
wire  signed [32:0] sext_ln813_298_fu_40816_p1;
wire  signed [32:0] sext_ln813_297_fu_40812_p1;
wire   [32:0] ret_V_157_fu_40820_p2;
wire   [31:0] p_Val2_799_fu_40834_p2;
wire   [0:0] p_Result_799_fu_40826_p3;
wire   [0:0] p_Result_800_fu_40840_p3;
wire   [0:0] xor_ln895_481_fu_40848_p2;
wire   [0:0] xor_ln896_481_fu_40860_p2;
wire   [0:0] xor_ln302_315_fu_40872_p2;
wire   [0:0] overflow_319_fu_40854_p2;
wire   [0:0] xor_ln302_316_fu_40878_p2;
wire   [0:0] underflow_319_fu_40866_p2;
wire   [0:0] or_ln302_157_fu_40884_p2;
wire   [31:0] select_ln302_315_fu_40890_p3;
wire   [31:0] select_ln350_157_fu_40898_p3;
wire  signed [31:0] lhs_140_fu_40094_p3;
wire  signed [31:0] rhs_158_fu_39228_p3;
wire  signed [32:0] sext_ln813_300_fu_40918_p1;
wire  signed [32:0] sext_ln813_299_fu_40914_p1;
wire   [32:0] ret_V_158_fu_40922_p2;
wire   [31:0] p_Val2_801_fu_40936_p2;
wire   [0:0] p_Result_801_fu_40928_p3;
wire   [0:0] p_Result_802_fu_40942_p3;
wire   [0:0] xor_ln895_482_fu_40950_p2;
wire   [0:0] xor_ln896_482_fu_40962_p2;
wire   [0:0] xor_ln302_317_fu_40974_p2;
wire   [0:0] overflow_320_fu_40956_p2;
wire   [0:0] xor_ln302_318_fu_40980_p2;
wire   [0:0] underflow_320_fu_40968_p2;
wire   [0:0] or_ln302_158_fu_40986_p2;
wire   [31:0] select_ln302_317_fu_40992_p3;
wire   [31:0] select_ln350_158_fu_41000_p3;
wire  signed [31:0] lhs_141_fu_40194_p3;
wire  signed [31:0] rhs_159_fu_39246_p3;
wire  signed [32:0] sext_ln813_302_fu_41020_p1;
wire  signed [32:0] sext_ln813_301_fu_41016_p1;
wire   [32:0] ret_V_159_fu_41024_p2;
wire   [31:0] p_Val2_803_fu_41038_p2;
wire   [0:0] p_Result_803_fu_41030_p3;
wire   [0:0] p_Result_804_fu_41044_p3;
wire   [0:0] xor_ln895_483_fu_41052_p2;
wire   [0:0] xor_ln896_483_fu_41064_p2;
wire   [0:0] xor_ln302_319_fu_41076_p2;
wire   [0:0] overflow_321_fu_41058_p2;
wire   [0:0] xor_ln302_320_fu_41082_p2;
wire   [0:0] underflow_321_fu_41070_p2;
wire   [0:0] or_ln302_159_fu_41088_p2;
wire   [31:0] select_ln302_319_fu_41094_p3;
wire   [31:0] select_ln350_159_fu_41102_p3;
wire  signed [31:0] lhs_142_fu_40294_p3;
wire  signed [31:0] rhs_160_fu_39394_p3;
wire  signed [32:0] sext_ln813_304_fu_41122_p1;
wire  signed [32:0] sext_ln813_303_fu_41118_p1;
wire   [32:0] ret_V_160_fu_41126_p2;
wire   [31:0] p_Val2_805_fu_41140_p2;
wire   [0:0] p_Result_805_fu_41132_p3;
wire   [0:0] p_Result_806_fu_41146_p3;
wire   [0:0] xor_ln895_484_fu_41154_p2;
wire   [0:0] xor_ln896_484_fu_41166_p2;
wire   [0:0] xor_ln302_321_fu_41178_p2;
wire   [0:0] overflow_322_fu_41160_p2;
wire   [0:0] xor_ln302_322_fu_41184_p2;
wire   [0:0] underflow_322_fu_41172_p2;
wire   [0:0] or_ln302_160_fu_41190_p2;
wire   [31:0] select_ln302_321_fu_41196_p3;
wire   [31:0] select_ln350_160_fu_41204_p3;
wire   [31:0] select_ln302_306_fu_40396_p3;
wire   [31:0] select_ln302_308_fu_40498_p3;
wire   [31:0] select_ln302_310_fu_40600_p3;
wire   [31:0] select_ln302_312_fu_40702_p3;
wire   [31:0] select_ln302_314_fu_40804_p3;
wire   [31:0] select_ln302_316_fu_40906_p3;
wire   [31:0] select_ln302_318_fu_41008_p3;
wire   [31:0] select_ln302_320_fu_41110_p3;
wire   [31:0] select_ln302_322_fu_41212_p3;
reg    ap_ce_reg;
reg  signed [31:0] p_read_int_reg;
reg  signed [31:0] p_read1_int_reg;
reg  signed [31:0] p_read2_int_reg;
reg   [31:0] p_read3_int_reg;
reg   [31:0] p_read4_int_reg;
reg   [31:0] p_read5_int_reg;
reg   [31:0] p_read6_int_reg;
reg   [31:0] p_read7_int_reg;
reg   [31:0] p_read8_int_reg;
reg   [31:0] ap_return_0_int_reg;
reg   [31:0] ap_return_1_int_reg;
reg   [31:0] ap_return_2_int_reg;
reg   [31:0] ap_return_3_int_reg;
reg   [31:0] ap_return_4_int_reg;
reg   [31:0] ap_return_5_int_reg;
reg   [31:0] ap_return_6_int_reg;
reg   [31:0] ap_return_7_int_reg;
reg   [31:0] ap_return_8_int_reg;

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U48(
    .din0(r_V_124_fu_462_p0),
    .din1(r_V_124_fu_462_p1),
    .dout(r_V_124_fu_462_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U49(
    .din0(r_V_107_fu_463_p0),
    .din1(r_V_107_fu_463_p1),
    .dout(r_V_107_fu_463_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U50(
    .din0(p_read_29_reg_41293_pp0_iter1_reg),
    .din1(r_V_137_fu_464_p1),
    .dout(r_V_137_fu_464_p2)
);

motorB_mul_32s_21s_52_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 21 ),
    .dout_WIDTH( 52 ))
mul_32s_21s_52_1_0_U51(
    .din0(p_read2_int_reg),
    .din1(r_V_99_fu_465_p1),
    .dout(r_V_99_fu_465_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U52(
    .din0(r_V_104_fu_466_p0),
    .din1(r_V_104_fu_466_p1),
    .dout(r_V_104_fu_466_p2)
);

motorB_mul_32s_18s_50_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 18 ),
    .dout_WIDTH( 50 ))
mul_32s_18s_50_1_0_U53(
    .din0(r_V_157_fu_467_p0),
    .din1(r_V_157_fu_467_p1),
    .dout(r_V_157_fu_467_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U54(
    .din0(r_V_115_fu_468_p0),
    .din1(r_V_115_fu_468_p1),
    .dout(r_V_115_fu_468_p2)
);

motorB_mul_32s_15s_47_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 47 ))
mul_32s_15s_47_1_0_U55(
    .din0(p_read2_int_reg),
    .din1(r_V_103_fu_469_p1),
    .dout(r_V_103_fu_469_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U56(
    .din0(p_read_31_reg_41314),
    .din1(r_V_118_fu_470_p1),
    .dout(r_V_118_fu_470_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U57(
    .din0(r_V_112_fu_471_p0),
    .din1(r_V_112_fu_471_p1),
    .dout(r_V_112_fu_471_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U58(
    .din0(r_V_123_fu_472_p0),
    .din1(r_V_123_fu_472_p1),
    .dout(r_V_123_fu_472_p2)
);

motorB_mul_32s_18s_50_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 18 ),
    .dout_WIDTH( 50 ))
mul_32s_18s_50_1_0_U59(
    .din0(r_V_153_fu_473_p0),
    .din1(r_V_153_fu_473_p1),
    .dout(r_V_153_fu_473_p2)
);

motorB_mul_32s_9ns_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9ns_41_1_0_U60(
    .din0(r_V_102_fu_474_p0),
    .din1(r_V_102_fu_474_p1),
    .dout(r_V_102_fu_474_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U61(
    .din0(p_read_31_reg_41314),
    .din1(r_V_114_fu_475_p1),
    .dout(r_V_114_fu_475_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U62(
    .din0(r_V_145_fu_476_p0),
    .din1(r_V_145_fu_476_p1),
    .dout(r_V_145_fu_476_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U63(
    .din0(r_V_121_fu_477_p0),
    .din1(r_V_121_fu_477_p1),
    .dout(r_V_121_fu_477_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U64(
    .din0(p_read2_int_reg),
    .din1(r_V_101_fu_478_p1),
    .dout(r_V_101_fu_478_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U65(
    .din0(r_V_127_fu_479_p0),
    .din1(r_V_127_fu_479_p1),
    .dout(r_V_127_fu_479_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U66(
    .din0(r_V_90_fu_480_p0),
    .din1(r_V_90_fu_480_p1),
    .dout(r_V_90_fu_480_p2)
);

motorB_mul_32s_24s_55_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 24 ),
    .dout_WIDTH( 55 ))
mul_32s_24s_55_1_0_U67(
    .din0(p_read_28_reg_41284_pp0_iter2_reg),
    .din1(r_V_140_fu_481_p1),
    .dout(r_V_140_fu_481_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U68(
    .din0(p_read1_int_reg),
    .din1(r_V_89_fu_482_p1),
    .dout(r_V_89_fu_482_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U69(
    .din0(r_V_155_fu_483_p0),
    .din1(r_V_155_fu_483_p1),
    .dout(r_V_155_fu_483_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U70(
    .din0(r_V_79_fu_484_p0),
    .din1(r_V_79_fu_484_p1),
    .dout(r_V_79_fu_484_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U71(
    .din0(r_V_109_fu_485_p0),
    .din1(r_V_109_fu_485_p1),
    .dout(r_V_109_fu_485_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U72(
    .din0(r_V_133_fu_486_p0),
    .din1(r_V_133_fu_486_p1),
    .dout(r_V_133_fu_486_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U73(
    .din0(r_V_81_fu_489_p0),
    .din1(r_V_81_fu_489_p1),
    .dout(r_V_81_fu_489_p2)
);

motorB_mul_32s_17ns_49_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 17 ),
    .dout_WIDTH( 49 ))
mul_32s_17ns_49_1_0_U74(
    .din0(r_V_144_fu_490_p0),
    .din1(r_V_144_fu_490_p1),
    .dout(r_V_144_fu_490_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U75(
    .din0(p_read_30_reg_41303_pp0_iter1_reg),
    .din1(r_V_130_fu_491_p1),
    .dout(r_V_130_fu_491_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U76(
    .din0(p_read_28_reg_41284_pp0_iter2_reg),
    .din1(r_V_142_fu_492_p1),
    .dout(r_V_142_fu_492_p2)
);

motorB_mul_32s_24ns_55_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 24 ),
    .dout_WIDTH( 55 ))
mul_32s_24ns_55_1_0_U77(
    .din0(p_read_27_reg_41274_pp0_iter2_reg),
    .din1(r_V_149_fu_493_p1),
    .dout(r_V_149_fu_493_p2)
);

motorB_mul_32s_8s_40_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 40 ))
mul_32s_8s_40_1_0_U78(
    .din0(p_read_int_reg),
    .din1(r_V_84_fu_494_p1),
    .dout(r_V_84_fu_494_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U79(
    .din0(r_V_85_fu_495_p0),
    .din1(r_V_85_fu_495_p1),
    .dout(r_V_85_fu_495_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U80(
    .din0(r_V_135_fu_496_p0),
    .din1(r_V_135_fu_496_p1),
    .dout(r_V_135_fu_496_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U81(
    .din0(r_V_82_fu_497_p0),
    .din1(r_V_82_fu_497_p1),
    .dout(r_V_82_fu_497_p2)
);

motorB_mul_32s_8s_40_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 40 ))
mul_32s_8s_40_1_0_U82(
    .din0(p_read1_int_reg),
    .din1(r_V_88_fu_498_p1),
    .dout(r_V_88_fu_498_p2)
);

motorB_mul_32s_7s_39_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 39 ))
mul_32s_7s_39_1_0_U83(
    .din0(p_read1_int_reg),
    .din1(r_V_94_fu_499_p1),
    .dout(r_V_94_fu_499_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U84(
    .din0(r_V_136_fu_500_p0),
    .din1(r_V_136_fu_500_p1),
    .dout(r_V_136_fu_500_p2)
);

motorB_mul_32s_25ns_56_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 25 ),
    .dout_WIDTH( 56 ))
mul_32s_25ns_56_1_0_U85(
    .din0(p_read2_int_reg),
    .din1(r_V_98_fu_501_p1),
    .dout(r_V_98_fu_501_p2)
);

motorB_mul_32s_24s_55_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 24 ),
    .dout_WIDTH( 55 ))
mul_32s_24s_55_1_0_U86(
    .din0(p_read2_int_reg),
    .din1(r_V_95_fu_503_p1),
    .dout(r_V_95_fu_503_p2)
);

motorB_mul_32s_9ns_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9ns_41_1_0_U87(
    .din0(r_V_97_fu_504_p0),
    .din1(r_V_97_fu_504_p1),
    .dout(r_V_97_fu_504_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U88(
    .din0(p_read1_int_reg),
    .din1(r_V_86_fu_505_p1),
    .dout(r_V_86_fu_505_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U89(
    .din0(r_V_131_fu_506_p0),
    .din1(r_V_131_fu_506_p1),
    .dout(r_V_131_fu_506_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U90(
    .din0(p_read_int_reg),
    .din1(r_V_83_fu_507_p1),
    .dout(r_V_83_fu_507_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U91(
    .din0(r_V_147_fu_508_p0),
    .din1(r_V_147_fu_508_p1),
    .dout(r_V_147_fu_508_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U92(
    .din0(r_V_80_fu_509_p0),
    .din1(r_V_80_fu_509_p1),
    .dout(r_V_80_fu_509_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U93(
    .din0(r_V_125_fu_510_p0),
    .din1(r_V_125_fu_510_p1),
    .dout(r_V_125_fu_510_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U94(
    .din0(r_V_106_fu_512_p0),
    .din1(r_V_106_fu_512_p1),
    .dout(r_V_106_fu_512_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U95(
    .din0(p_read_30_reg_41303_pp0_iter1_reg),
    .din1(r_V_128_fu_513_p1),
    .dout(r_V_128_fu_513_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U96(
    .din0(r_V_146_fu_514_p0),
    .din1(r_V_146_fu_514_p1),
    .dout(r_V_146_fu_514_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U97(
    .din0(r_V_126_fu_515_p0),
    .din1(r_V_126_fu_515_p1),
    .dout(r_V_126_fu_515_p2)
);

motorB_mul_32s_18ns_50_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 18 ),
    .dout_WIDTH( 50 ))
mul_32s_18ns_50_1_0_U98(
    .din0(r_V_152_fu_516_p0),
    .din1(r_V_152_fu_516_p1),
    .dout(r_V_152_fu_516_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U99(
    .din0(r_V_151_fu_517_p0),
    .din1(r_V_151_fu_517_p1),
    .dout(r_V_151_fu_517_p2)
);

motorB_mul_32s_17ns_49_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 17 ),
    .dout_WIDTH( 49 ))
mul_32s_17ns_49_1_0_U100(
    .din0(r_V_148_fu_518_p0),
    .din1(r_V_148_fu_518_p1),
    .dout(r_V_148_fu_518_p2)
);

motorB_mul_32s_15s_47_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 47 ))
mul_32s_15s_47_1_0_U101(
    .din0(p_read_31_reg_41314),
    .din1(r_V_117_fu_519_p1),
    .dout(r_V_117_fu_519_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U102(
    .din0(r_V_120_fu_520_p0),
    .din1(r_V_120_fu_520_p1),
    .dout(r_V_120_fu_520_p2)
);

motorB_mul_32s_8ns_40_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 40 ))
mul_32s_8ns_40_1_0_U103(
    .din0(p_read_30_reg_41303_pp0_iter1_reg),
    .din1(r_V_129_fu_521_p1),
    .dout(r_V_129_fu_521_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U104(
    .din0(r_V_92_fu_522_p0),
    .din1(r_V_92_fu_522_p1),
    .dout(r_V_92_fu_522_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U105(
    .din0(r_V_154_fu_523_p0),
    .din1(r_V_154_fu_523_p1),
    .dout(r_V_154_fu_523_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U106(
    .din0(r_V_134_fu_525_p0),
    .din1(r_V_134_fu_525_p1),
    .dout(r_V_134_fu_525_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U107(
    .din0(r_V_111_fu_526_p0),
    .din1(r_V_111_fu_526_p1),
    .dout(r_V_111_fu_526_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U108(
    .din0(r_V_78_fu_527_p0),
    .din1(r_V_78_fu_527_p1),
    .dout(r_V_78_fu_527_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U109(
    .din0(p_read_29_reg_41293_pp0_iter1_reg),
    .din1(r_V_138_fu_528_p1),
    .dout(r_V_138_fu_528_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U110(
    .din0(r_V_108_fu_529_p0),
    .din1(r_V_108_fu_529_p1),
    .dout(r_V_108_fu_529_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U111(
    .din0(p_read2_int_reg),
    .din1(r_V_96_fu_530_p1),
    .dout(r_V_96_fu_530_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U112(
    .din0(r_V_150_fu_531_p0),
    .din1(r_V_150_fu_531_p1),
    .dout(r_V_150_fu_531_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U113(
    .din0(p_read1_int_reg),
    .din1(r_V_93_fu_532_p1),
    .dout(r_V_93_fu_532_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U114(
    .din0(r_V_132_fu_533_p0),
    .din1(r_V_132_fu_533_p1),
    .dout(r_V_132_fu_533_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U115(
    .din0(p_read2_int_reg),
    .din1(r_V_100_fu_534_p1),
    .dout(r_V_100_fu_534_p2)
);

motorB_mul_32s_24ns_55_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 24 ),
    .dout_WIDTH( 55 ))
mul_32s_24ns_55_1_0_U116(
    .din0(p_read_31_reg_41314),
    .din1(r_V_113_fu_535_p1),
    .dout(r_V_113_fu_535_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U117(
    .din0(r_V_fu_536_p0),
    .din1(r_V_fu_536_p1),
    .dout(r_V_fu_536_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U118(
    .din0(r_V_116_fu_537_p0),
    .din1(r_V_116_fu_537_p1),
    .dout(r_V_116_fu_537_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U119(
    .din0(r_V_87_fu_538_p0),
    .din1(r_V_87_fu_538_p1),
    .dout(r_V_87_fu_538_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U120(
    .din0(r_V_105_fu_539_p0),
    .din1(r_V_105_fu_539_p1),
    .dout(r_V_105_fu_539_p2)
);

motorB_mul_32s_18s_50_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 18 ),
    .dout_WIDTH( 50 ))
mul_32s_18s_50_1_0_U121(
    .din0(p_read_28_reg_41284_pp0_iter2_reg),
    .din1(r_V_143_fu_540_p1),
    .dout(r_V_143_fu_540_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U122(
    .din0(r_V_141_fu_541_p0),
    .din1(r_V_141_fu_541_p1),
    .dout(r_V_141_fu_541_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U123(
    .din0(r_V_119_fu_542_p0),
    .din1(r_V_119_fu_542_p1),
    .dout(r_V_119_fu_542_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        Range2_all_ones_100_reg_41997 <= r_V_99_fu_465_p2[32'd51];
        Range2_all_ones_101_reg_42026 <= r_V_100_fu_534_p2[32'd44];
        Range2_all_ones_102_reg_42055 <= r_V_101_fu_478_p2[32'd42];
        Range2_all_ones_103_reg_42084 <= r_V_102_fu_474_p2[32'd40];
        Range2_all_ones_104_reg_42113 <= r_V_103_fu_469_p2[32'd46];
        Range2_all_ones_105_reg_42276 <= r_V_104_fu_466_p2[32'd41];
        Range2_all_ones_106_reg_42307 <= r_V_105_fu_539_p2[32'd42];
        Range2_all_ones_107_reg_42338 <= r_V_106_fu_512_p2[32'd41];
        Range2_all_ones_108_reg_42369 <= r_V_107_fu_463_p2[32'd42];
        Range2_all_ones_109_reg_42400 <= r_V_108_fu_529_p2[32'd43];
        Range2_all_ones_110_reg_42431 <= r_V_109_fu_485_p2[32'd41];
        Range2_all_ones_112_reg_42477 <= r_V_111_fu_526_p2[32'd43];
        Range2_all_ones_113_reg_42508 <= r_V_112_fu_471_p2[32'd42];
        Range2_all_ones_114_reg_42537 <= r_V_113_fu_535_p2[32'd54];
        Range2_all_ones_115_reg_42566 <= r_V_114_fu_475_p2[32'd41];
        Range2_all_ones_116_reg_42595 <= r_V_115_fu_468_p2[32'd44];
        Range2_all_ones_117_reg_42624 <= r_V_116_fu_537_p2[32'd44];
        Range2_all_ones_118_reg_42653 <= r_V_117_fu_519_p2[32'd46];
        Range2_all_ones_119_reg_42682 <= r_V_118_fu_470_p2[32'd42];
        Range2_all_ones_120_reg_42711 <= r_V_119_fu_542_p2[32'd44];
        Range2_all_ones_121_reg_42740 <= r_V_120_fu_520_p2[32'd43];
        Range2_all_ones_122_reg_42769 <= r_V_121_fu_477_p2[32'd43];
        Range2_all_ones_124_reg_42869 <= r_V_123_fu_472_p2[32'd42];
        Range2_all_ones_125_reg_42900 <= r_V_124_fu_462_p2[32'd43];
        Range2_all_ones_126_reg_42931 <= r_V_125_fu_510_p2[32'd42];
        Range2_all_ones_127_reg_42962 <= r_V_126_fu_515_p2[32'd43];
        Range2_all_ones_128_reg_42993 <= r_V_127_fu_479_p2[32'd42];
        Range2_all_ones_129_reg_43024 <= r_V_128_fu_513_p2[32'd44];
        Range2_all_ones_130_reg_43055 <= r_V_129_fu_521_p2[32'd39];
        Range2_all_ones_131_reg_43086 <= r_V_130_fu_491_p2[32'd41];
        Range2_all_ones_132_reg_43115 <= r_V_131_fu_506_p2[32'd43];
        Range2_all_ones_133_reg_43144 <= r_V_132_fu_533_p2[32'd42];
        Range2_all_ones_134_reg_43173 <= r_V_133_fu_486_p2[32'd42];
        Range2_all_ones_135_reg_43202 <= r_V_134_fu_525_p2[32'd43];
        Range2_all_ones_136_reg_43231 <= r_V_135_fu_496_p2[32'd42];
        Range2_all_ones_137_reg_43260 <= r_V_136_fu_500_p2[32'd42];
        Range2_all_ones_138_reg_43289 <= r_V_137_fu_464_p2[32'd40];
        Range2_all_ones_139_reg_43318 <= r_V_138_fu_528_p2[32'd41];
        Range2_all_ones_141_reg_43544 <= r_V_140_fu_481_p2[32'd54];
        Range2_all_ones_142_reg_43575 <= r_V_141_fu_541_p2[32'd43];
        Range2_all_ones_143_reg_43606 <= r_V_142_fu_492_p2[32'd42];
        Range2_all_ones_144_reg_43637 <= r_V_143_fu_540_p2[32'd49];
        Range2_all_ones_145_reg_43668 <= r_V_144_fu_490_p2[32'd48];
        Range2_all_ones_146_reg_43699 <= r_V_145_fu_476_p2[32'd43];
        Range2_all_ones_147_reg_43730 <= r_V_146_fu_514_p2[32'd43];
        Range2_all_ones_148_reg_43761 <= r_V_147_fu_508_p2[32'd43];
        Range2_all_ones_149_reg_43792 <= r_V_148_fu_518_p2[32'd48];
        Range2_all_ones_150_reg_43821 <= r_V_149_fu_493_p2[32'd54];
        Range2_all_ones_151_reg_43850 <= r_V_150_fu_531_p2[32'd41];
        Range2_all_ones_152_reg_43879 <= r_V_151_fu_517_p2[32'd43];
        Range2_all_ones_153_reg_43908 <= r_V_152_fu_516_p2[32'd49];
        Range2_all_ones_154_reg_43937 <= r_V_153_fu_473_p2[32'd49];
        Range2_all_ones_155_reg_43966 <= r_V_154_fu_523_p2[32'd41];
        Range2_all_ones_156_reg_43995 <= r_V_155_fu_483_p2[32'd43];
        Range2_all_ones_158_reg_44039 <= r_V_157_fu_467_p2[32'd49];
        Range2_all_ones_79_reg_41388 <= r_V_78_fu_527_p2[32'd42];
        Range2_all_ones_80_reg_41419 <= r_V_79_fu_484_p2[32'd43];
        Range2_all_ones_81_reg_41450 <= r_V_80_fu_509_p2[32'd41];
        Range2_all_ones_82_reg_41481 <= r_V_81_fu_489_p2[32'd41];
        Range2_all_ones_83_reg_41512 <= r_V_82_fu_497_p2[32'd43];
        Range2_all_ones_84_reg_41543 <= r_V_83_fu_507_p2[32'd44];
        Range2_all_ones_85_reg_41574 <= r_V_84_fu_494_p2[32'd39];
        Range2_all_ones_86_reg_41605 <= r_V_85_fu_495_p2[32'd42];
        Range2_all_ones_87_reg_41634 <= r_V_86_fu_505_p2[32'd44];
        Range2_all_ones_88_reg_41663 <= r_V_87_fu_538_p2[32'd41];
        Range2_all_ones_89_reg_41692 <= r_V_88_fu_498_p2[32'd39];
        Range2_all_ones_90_reg_41721 <= r_V_89_fu_482_p2[32'd43];
        Range2_all_ones_91_reg_41750 <= r_V_90_fu_480_p2[32'd41];
        Range2_all_ones_93_reg_41794 <= r_V_92_fu_522_p2[32'd41];
        Range2_all_ones_94_reg_41823 <= r_V_93_fu_532_p2[32'd42];
        Range2_all_ones_95_reg_41852 <= r_V_94_fu_499_p2[32'd38];
        Range2_all_ones_96_reg_41881 <= r_V_95_fu_503_p2[32'd54];
        Range2_all_ones_97_reg_41910 <= r_V_96_fu_530_p2[32'd43];
        Range2_all_ones_98_reg_41939 <= r_V_97_fu_504_p2[32'd40];
        Range2_all_ones_99_reg_41968 <= r_V_98_fu_501_p2[32'd55];
        Range2_all_ones_reg_41357 <= r_V_fu_536_p2[32'd41];
        lhs_125_reg_44046 <= lhs_125_fu_36252_p3;
        lhs_126_reg_44052 <= lhs_126_fu_36354_p3;
        lhs_127_reg_44058 <= lhs_127_fu_36456_p3;
        lhs_128_reg_44064 <= lhs_128_fu_36558_p3;
        lhs_129_reg_44070 <= lhs_129_fu_36660_p3;
        lhs_130_reg_44076 <= lhs_130_fu_36762_p3;
        lhs_131_reg_44082 <= lhs_131_fu_36864_p3;
        lhs_132_reg_44088 <= lhs_132_fu_36966_p3;
        lhs_133_reg_44094 <= lhs_133_fu_37068_p3;
        lhs_80_reg_42776 <= lhs_80_fu_24598_p3;
        lhs_81_reg_42782 <= lhs_81_fu_24700_p3;
        lhs_82_reg_42788 <= lhs_82_fu_24802_p3;
        lhs_83_reg_42794 <= lhs_83_fu_24904_p3;
        lhs_84_reg_42800 <= lhs_84_fu_25006_p3;
        lhs_85_reg_42806 <= lhs_85_fu_25108_p3;
        lhs_86_reg_42812 <= lhs_86_fu_25210_p3;
        lhs_87_reg_42818 <= lhs_87_fu_25312_p3;
        lhs_88_reg_42824 <= lhs_88_fu_25414_p3;
        or_ln346_100_reg_42166 <= or_ln346_100_fu_21697_p2;
        or_ln346_102_reg_42187 <= or_ln346_102_fu_21967_p2;
        or_ln346_103_reg_42202 <= or_ln346_103_fu_22096_p2;
        or_ln346_104_reg_42217 <= or_ln346_104_fu_22225_p2;
        or_ln346_105_reg_42232 <= or_ln346_105_fu_22354_p2;
        or_ln346_106_reg_42247 <= or_ln346_106_fu_22483_p2;
        or_ln346_113_reg_42448 <= or_ln346_113_fu_23083_p2;
        or_ln346_125_reg_42840 <= or_ln346_125_fu_28111_p2;
        or_ln346_142_reg_43335 <= or_ln346_142_fu_29178_p2;
        or_ln346_159_reg_44012 <= or_ln346_159_fu_34670_p2;
        or_ln346_94_reg_41767 <= or_ln346_94_fu_18301_p2;
        or_ln346_99_reg_42151 <= or_ln346_99_fu_21568_p2;
        overflow_175_reg_41762 <= overflow_175_fu_18271_p2;
        overflow_180_reg_42146 <= overflow_180_fu_21539_p2;
        overflow_181_reg_42161 <= overflow_181_fu_21668_p2;
        overflow_183_reg_42182 <= overflow_183_fu_21938_p2;
        overflow_184_reg_42197 <= overflow_184_fu_22067_p2;
        overflow_185_reg_42212 <= overflow_185_fu_22196_p2;
        overflow_186_reg_42227 <= overflow_186_fu_22325_p2;
        overflow_187_reg_42242 <= overflow_187_fu_22454_p2;
        overflow_194_reg_42443 <= overflow_194_fu_23053_p2;
        overflow_206_reg_42835 <= overflow_206_fu_28081_p2;
        overflow_223_reg_43330 <= overflow_223_fu_29148_p2;
        overflow_240_reg_44007 <= overflow_240_fu_34640_p2;
        p_Result_403_reg_41339 <= r_V_fu_536_p2[32'd41];
        p_Result_404_reg_41350 <= p_Val2_403_fu_17315_p2[32'd18];
        p_Result_405_reg_41364 <= r_V_78_fu_527_p2[32'd42];
        p_Result_406_reg_41370 <= r_V_78_fu_527_p2[32'd42];
        p_Result_407_reg_41381 <= p_Val2_406_fu_17379_p2[32'd19];
        p_Result_408_reg_41395 <= r_V_79_fu_484_p2[32'd43];
        p_Result_409_reg_41401 <= r_V_79_fu_484_p2[32'd43];
        p_Result_410_reg_41412 <= p_Val2_409_fu_17443_p2[32'd20];
        p_Result_411_reg_41426 <= r_V_80_fu_509_p2[32'd41];
        p_Result_412_reg_41432 <= r_V_80_fu_509_p2[32'd41];
        p_Result_413_reg_41443 <= p_Val2_412_fu_17507_p2[32'd18];
        p_Result_414_reg_41457 <= r_V_81_fu_489_p2[32'd41];
        p_Result_415_reg_41463 <= r_V_81_fu_489_p2[32'd41];
        p_Result_416_reg_41474 <= p_Val2_415_fu_17571_p2[32'd18];
        p_Result_417_reg_41488 <= r_V_82_fu_497_p2[32'd43];
        p_Result_418_reg_41494 <= r_V_82_fu_497_p2[32'd43];
        p_Result_419_reg_41505 <= p_Val2_418_fu_17635_p2[32'd20];
        p_Result_420_reg_41519 <= r_V_83_fu_507_p2[32'd44];
        p_Result_421_reg_41525 <= r_V_83_fu_507_p2[32'd44];
        p_Result_422_reg_41536 <= p_Val2_421_fu_17699_p2[32'd21];
        p_Result_423_reg_41550 <= r_V_84_fu_494_p2[32'd39];
        p_Result_424_reg_41556 <= r_V_84_fu_494_p2[32'd39];
        p_Result_425_reg_41567 <= p_Val2_424_fu_17763_p2[32'd16];
        p_Result_426_reg_41581 <= r_V_85_fu_495_p2[32'd42];
        p_Result_427_reg_41587 <= r_V_85_fu_495_p2[32'd42];
        p_Result_428_reg_41598 <= p_Val2_427_fu_17827_p2[32'd19];
        p_Result_429_reg_41612 <= r_V_86_fu_505_p2[32'd44];
        p_Result_430_reg_41623 <= r_V_86_fu_505_p2[32'd44];
        p_Result_432_reg_41641 <= r_V_87_fu_538_p2[32'd41];
        p_Result_433_reg_41652 <= r_V_87_fu_538_p2[32'd41];
        p_Result_435_reg_41670 <= r_V_88_fu_498_p2[32'd39];
        p_Result_436_reg_41681 <= r_V_88_fu_498_p2[32'd39];
        p_Result_438_reg_41699 <= r_V_89_fu_482_p2[32'd43];
        p_Result_439_reg_41710 <= r_V_89_fu_482_p2[32'd43];
        p_Result_441_reg_41728 <= r_V_90_fu_480_p2[32'd41];
        p_Result_442_reg_41739 <= r_V_90_fu_480_p2[32'd41];
        p_Result_447_reg_41772 <= r_V_92_fu_522_p2[32'd41];
        p_Result_448_reg_41783 <= r_V_92_fu_522_p2[32'd41];
        p_Result_450_reg_41801 <= r_V_93_fu_532_p2[32'd42];
        p_Result_451_reg_41812 <= r_V_93_fu_532_p2[32'd42];
        p_Result_453_reg_41830 <= r_V_94_fu_499_p2[32'd38];
        p_Result_454_reg_41841 <= r_V_94_fu_499_p2[32'd38];
        p_Result_456_reg_41859 <= r_V_95_fu_503_p2[32'd54];
        p_Result_457_reg_41870 <= r_V_95_fu_503_p2[32'd54];
        p_Result_459_reg_41888 <= r_V_96_fu_530_p2[32'd43];
        p_Result_460_reg_41899 <= r_V_96_fu_530_p2[32'd43];
        p_Result_462_reg_41917 <= r_V_97_fu_504_p2[32'd40];
        p_Result_463_reg_41928 <= r_V_97_fu_504_p2[32'd40];
        p_Result_465_reg_41946 <= r_V_98_fu_501_p2[32'd55];
        p_Result_466_reg_41957 <= r_V_98_fu_501_p2[32'd55];
        p_Result_468_reg_41975 <= r_V_99_fu_465_p2[32'd51];
        p_Result_469_reg_41986 <= r_V_99_fu_465_p2[32'd51];
        p_Result_471_reg_42004 <= r_V_100_fu_534_p2[32'd44];
        p_Result_472_reg_42015 <= r_V_100_fu_534_p2[32'd44];
        p_Result_474_reg_42033 <= r_V_101_fu_478_p2[32'd42];
        p_Result_475_reg_42044 <= r_V_101_fu_478_p2[32'd42];
        p_Result_477_reg_42062 <= r_V_102_fu_474_p2[32'd40];
        p_Result_478_reg_42073 <= r_V_102_fu_474_p2[32'd40];
        p_Result_480_reg_42091 <= r_V_103_fu_469_p2[32'd46];
        p_Result_481_reg_42102 <= r_V_103_fu_469_p2[32'd46];
        p_Result_483_reg_42252 <= r_V_104_fu_466_p2[32'd41];
        p_Result_484_reg_42258 <= r_V_104_fu_466_p2[32'd41];
        p_Result_485_reg_42269 <= p_Val2_484_fu_22548_p2[32'd18];
        p_Result_486_reg_42283 <= r_V_105_fu_539_p2[32'd42];
        p_Result_487_reg_42289 <= r_V_105_fu_539_p2[32'd42];
        p_Result_488_reg_42300 <= p_Val2_487_fu_22612_p2[32'd19];
        p_Result_489_reg_42314 <= r_V_106_fu_512_p2[32'd41];
        p_Result_490_reg_42320 <= r_V_106_fu_512_p2[32'd41];
        p_Result_491_reg_42331 <= p_Val2_490_fu_22676_p2[32'd18];
        p_Result_492_reg_42345 <= r_V_107_fu_463_p2[32'd42];
        p_Result_493_reg_42351 <= r_V_107_fu_463_p2[32'd42];
        p_Result_494_reg_42362 <= p_Val2_493_fu_22740_p2[32'd19];
        p_Result_495_reg_42376 <= r_V_108_fu_529_p2[32'd43];
        p_Result_496_reg_42382 <= r_V_108_fu_529_p2[32'd43];
        p_Result_497_reg_42393 <= p_Val2_496_fu_22804_p2[32'd20];
        p_Result_498_reg_42407 <= r_V_109_fu_485_p2[32'd41];
        p_Result_499_reg_42413 <= r_V_109_fu_485_p2[32'd41];
        p_Result_500_reg_42424 <= p_Val2_499_fu_22868_p2[32'd18];
        p_Result_504_reg_42453 <= r_V_111_fu_526_p2[32'd43];
        p_Result_505_reg_42459 <= r_V_111_fu_526_p2[32'd43];
        p_Result_506_reg_42470 <= p_Val2_505_fu_23131_p2[32'd20];
        p_Result_507_reg_42484 <= r_V_112_fu_471_p2[32'd42];
        p_Result_508_reg_42490 <= r_V_112_fu_471_p2[32'd42];
        p_Result_509_reg_42501 <= p_Val2_508_fu_23195_p2[32'd19];
        p_Result_510_reg_42515 <= r_V_113_fu_535_p2[32'd54];
        p_Result_511_reg_42526 <= r_V_113_fu_535_p2[32'd54];
        p_Result_513_reg_42544 <= r_V_114_fu_475_p2[32'd41];
        p_Result_514_reg_42555 <= r_V_114_fu_475_p2[32'd41];
        p_Result_516_reg_42573 <= r_V_115_fu_468_p2[32'd44];
        p_Result_517_reg_42584 <= r_V_115_fu_468_p2[32'd44];
        p_Result_519_reg_42602 <= r_V_116_fu_537_p2[32'd44];
        p_Result_520_reg_42613 <= r_V_116_fu_537_p2[32'd44];
        p_Result_522_reg_42631 <= r_V_117_fu_519_p2[32'd46];
        p_Result_523_reg_42642 <= r_V_117_fu_519_p2[32'd46];
        p_Result_525_reg_42660 <= r_V_118_fu_470_p2[32'd42];
        p_Result_526_reg_42671 <= r_V_118_fu_470_p2[32'd42];
        p_Result_528_reg_42689 <= r_V_119_fu_542_p2[32'd44];
        p_Result_529_reg_42700 <= r_V_119_fu_542_p2[32'd44];
        p_Result_531_reg_42718 <= r_V_120_fu_520_p2[32'd43];
        p_Result_532_reg_42729 <= r_V_120_fu_520_p2[32'd43];
        p_Result_534_reg_42747 <= r_V_121_fu_477_p2[32'd43];
        p_Result_535_reg_42758 <= r_V_121_fu_477_p2[32'd43];
        p_Result_540_reg_42845 <= r_V_123_fu_472_p2[32'd42];
        p_Result_541_reg_42851 <= r_V_123_fu_472_p2[32'd42];
        p_Result_542_reg_42862 <= p_Val2_541_fu_28159_p2[32'd19];
        p_Result_543_reg_42876 <= r_V_124_fu_462_p2[32'd43];
        p_Result_544_reg_42882 <= r_V_124_fu_462_p2[32'd43];
        p_Result_545_reg_42893 <= p_Val2_544_fu_28223_p2[32'd20];
        p_Result_546_reg_42907 <= r_V_125_fu_510_p2[32'd42];
        p_Result_547_reg_42913 <= r_V_125_fu_510_p2[32'd42];
        p_Result_548_reg_42924 <= p_Val2_547_fu_28287_p2[32'd19];
        p_Result_549_reg_42938 <= r_V_126_fu_515_p2[32'd43];
        p_Result_550_reg_42944 <= r_V_126_fu_515_p2[32'd43];
        p_Result_551_reg_42955 <= p_Val2_550_fu_28351_p2[32'd20];
        p_Result_552_reg_42969 <= r_V_127_fu_479_p2[32'd42];
        p_Result_553_reg_42975 <= r_V_127_fu_479_p2[32'd42];
        p_Result_554_reg_42986 <= p_Val2_553_fu_28415_p2[32'd19];
        p_Result_555_reg_43000 <= r_V_128_fu_513_p2[32'd44];
        p_Result_556_reg_43006 <= r_V_128_fu_513_p2[32'd44];
        p_Result_557_reg_43017 <= p_Val2_556_fu_28479_p2[32'd21];
        p_Result_558_reg_43031 <= r_V_129_fu_521_p2[32'd39];
        p_Result_559_reg_43037 <= r_V_129_fu_521_p2[32'd39];
        p_Result_560_reg_43048 <= p_Val2_559_fu_28543_p2[32'd16];
        p_Result_561_reg_43062 <= r_V_130_fu_491_p2[32'd41];
        p_Result_562_reg_43068 <= r_V_130_fu_491_p2[32'd41];
        p_Result_563_reg_43079 <= p_Val2_562_fu_28607_p2[32'd18];
        p_Result_564_reg_43093 <= r_V_131_fu_506_p2[32'd43];
        p_Result_565_reg_43104 <= r_V_131_fu_506_p2[32'd43];
        p_Result_567_reg_43122 <= r_V_132_fu_533_p2[32'd42];
        p_Result_568_reg_43133 <= r_V_132_fu_533_p2[32'd42];
        p_Result_570_reg_43151 <= r_V_133_fu_486_p2[32'd42];
        p_Result_571_reg_43162 <= r_V_133_fu_486_p2[32'd42];
        p_Result_573_reg_43180 <= r_V_134_fu_525_p2[32'd43];
        p_Result_574_reg_43191 <= r_V_134_fu_525_p2[32'd43];
        p_Result_576_reg_43209 <= r_V_135_fu_496_p2[32'd42];
        p_Result_577_reg_43220 <= r_V_135_fu_496_p2[32'd42];
        p_Result_579_reg_43238 <= r_V_136_fu_500_p2[32'd42];
        p_Result_580_reg_43249 <= r_V_136_fu_500_p2[32'd42];
        p_Result_582_reg_43267 <= r_V_137_fu_464_p2[32'd40];
        p_Result_583_reg_43278 <= r_V_137_fu_464_p2[32'd40];
        p_Result_585_reg_43296 <= r_V_138_fu_528_p2[32'd41];
        p_Result_586_reg_43307 <= r_V_138_fu_528_p2[32'd41];
        p_Result_591_reg_43520 <= r_V_140_fu_481_p2[32'd54];
        p_Result_592_reg_43526 <= r_V_140_fu_481_p2[32'd54];
        p_Result_593_reg_43537 <= p_Val2_592_fu_33614_p2[32'd31];
        p_Result_594_reg_43551 <= r_V_141_fu_541_p2[32'd43];
        p_Result_595_reg_43557 <= r_V_141_fu_541_p2[32'd43];
        p_Result_596_reg_43568 <= p_Val2_595_fu_33678_p2[32'd20];
        p_Result_597_reg_43582 <= r_V_142_fu_492_p2[32'd42];
        p_Result_598_reg_43588 <= r_V_142_fu_492_p2[32'd42];
        p_Result_599_reg_43599 <= p_Val2_598_fu_33742_p2[32'd19];
        p_Result_600_reg_43613 <= r_V_143_fu_540_p2[32'd49];
        p_Result_601_reg_43619 <= r_V_143_fu_540_p2[32'd49];
        p_Result_602_reg_43630 <= p_Val2_601_fu_33806_p2[32'd26];
        p_Result_603_reg_43644 <= r_V_144_fu_490_p2[32'd48];
        p_Result_604_reg_43650 <= r_V_144_fu_490_p2[32'd48];
        p_Result_605_reg_43661 <= p_Val2_604_fu_33870_p2[32'd25];
        p_Result_606_reg_43675 <= r_V_145_fu_476_p2[32'd43];
        p_Result_607_reg_43681 <= r_V_145_fu_476_p2[32'd43];
        p_Result_608_reg_43692 <= p_Val2_607_fu_33934_p2[32'd20];
        p_Result_609_reg_43706 <= r_V_146_fu_514_p2[32'd43];
        p_Result_610_reg_43712 <= r_V_146_fu_514_p2[32'd43];
        p_Result_611_reg_43723 <= p_Val2_610_fu_33998_p2[32'd20];
        p_Result_612_reg_43737 <= r_V_147_fu_508_p2[32'd43];
        p_Result_613_reg_43743 <= r_V_147_fu_508_p2[32'd43];
        p_Result_614_reg_43754 <= p_Val2_613_fu_34062_p2[32'd20];
        p_Result_615_reg_43768 <= r_V_148_fu_518_p2[32'd48];
        p_Result_616_reg_43774 <= r_V_148_fu_518_p2[32'd48];
        p_Result_617_reg_43785 <= p_Val2_616_fu_34126_p2[32'd25];
        p_Result_618_reg_43799 <= r_V_149_fu_493_p2[32'd54];
        p_Result_619_reg_43810 <= r_V_149_fu_493_p2[32'd54];
        p_Result_621_reg_43828 <= r_V_150_fu_531_p2[32'd41];
        p_Result_622_reg_43839 <= r_V_150_fu_531_p2[32'd41];
        p_Result_624_reg_43857 <= r_V_151_fu_517_p2[32'd43];
        p_Result_625_reg_43868 <= r_V_151_fu_517_p2[32'd43];
        p_Result_627_reg_43886 <= r_V_152_fu_516_p2[32'd49];
        p_Result_628_reg_43897 <= r_V_152_fu_516_p2[32'd49];
        p_Result_630_reg_43915 <= r_V_153_fu_473_p2[32'd49];
        p_Result_631_reg_43926 <= r_V_153_fu_473_p2[32'd49];
        p_Result_633_reg_43944 <= r_V_154_fu_523_p2[32'd41];
        p_Result_634_reg_43955 <= r_V_154_fu_523_p2[32'd41];
        p_Result_636_reg_43973 <= r_V_155_fu_483_p2[32'd43];
        p_Result_637_reg_43984 <= r_V_155_fu_483_p2[32'd43];
        p_Result_642_reg_44017 <= r_V_157_fu_467_p2[32'd49];
        p_Result_643_reg_44028 <= r_V_157_fu_467_p2[32'd49];
        p_Result_717_reg_43340 <= ret_V_116_fu_31006_p2[32'd32];
        p_Result_718_reg_43353 <= p_Val2_717_fu_31020_p2[32'd31];
        p_Result_719_reg_43360 <= ret_V_117_fu_31042_p2[32'd32];
        p_Result_720_reg_43373 <= p_Val2_719_fu_31056_p2[32'd31];
        p_Result_721_reg_43380 <= ret_V_118_fu_31078_p2[32'd32];
        p_Result_722_reg_43393 <= p_Val2_721_fu_31092_p2[32'd31];
        p_Result_723_reg_43400 <= ret_V_119_fu_31114_p2[32'd32];
        p_Result_724_reg_43413 <= p_Val2_723_fu_31128_p2[32'd31];
        p_Result_725_reg_43420 <= ret_V_120_fu_31150_p2[32'd32];
        p_Result_726_reg_43433 <= p_Val2_725_fu_31164_p2[32'd31];
        p_Result_727_reg_43440 <= ret_V_121_fu_31186_p2[32'd32];
        p_Result_728_reg_43453 <= p_Val2_727_fu_31200_p2[32'd31];
        p_Result_729_reg_43460 <= ret_V_122_fu_31222_p2[32'd32];
        p_Result_730_reg_43473 <= p_Val2_729_fu_31236_p2[32'd31];
        p_Result_731_reg_43480 <= ret_V_123_fu_31258_p2[32'd32];
        p_Result_732_reg_43493 <= p_Val2_731_fu_31272_p2[32'd31];
        p_Result_733_reg_43500 <= ret_V_124_fu_31294_p2[32'd32];
        p_Result_734_reg_43513 <= p_Val2_733_fu_31308_p2[32'd31];
        p_Result_s_reg_41333 <= r_V_fu_536_p2[32'd41];
        p_Val2_403_reg_41345 <= p_Val2_403_fu_17315_p2;
        p_Val2_406_reg_41376 <= p_Val2_406_fu_17379_p2;
        p_Val2_409_reg_41407 <= p_Val2_409_fu_17443_p2;
        p_Val2_412_reg_41438 <= p_Val2_412_fu_17507_p2;
        p_Val2_415_reg_41469 <= p_Val2_415_fu_17571_p2;
        p_Val2_418_reg_41500 <= p_Val2_418_fu_17635_p2;
        p_Val2_421_reg_41531 <= p_Val2_421_fu_17699_p2;
        p_Val2_424_reg_41562 <= p_Val2_424_fu_17763_p2;
        p_Val2_427_reg_41593 <= p_Val2_427_fu_17827_p2;
        p_Val2_429_reg_41618 <= {{r_V_86_fu_505_p2[44:24]}};
        p_Val2_432_reg_41647 <= {{r_V_87_fu_538_p2[41:24]}};
        p_Val2_435_reg_41676 <= {{r_V_88_fu_498_p2[39:24]}};
        p_Val2_438_reg_41705 <= {{r_V_89_fu_482_p2[43:24]}};
        p_Val2_441_reg_41734 <= {{r_V_90_fu_480_p2[41:24]}};
        p_Val2_445_reg_41757 <= p_Val2_445_fu_18169_p2;
        p_Val2_447_reg_41778 <= {{r_V_92_fu_522_p2[41:24]}};
        p_Val2_450_reg_41807 <= {{r_V_93_fu_532_p2[42:24]}};
        p_Val2_453_reg_41836 <= {{r_V_94_fu_499_p2[38:24]}};
        p_Val2_456_reg_41865 <= {{r_V_95_fu_503_p2[54:24]}};
        p_Val2_459_reg_41894 <= {{r_V_96_fu_530_p2[43:24]}};
        p_Val2_460_reg_42141 <= p_Val2_460_fu_21451_p2;
        p_Val2_462_reg_41923 <= {{r_V_97_fu_504_p2[40:24]}};
        p_Val2_463_reg_42156 <= p_Val2_463_fu_21580_p2;
        p_Val2_465_reg_41952 <= {{r_V_98_fu_501_p2[55:24]}};
        p_Val2_468_reg_41981 <= {{r_V_99_fu_465_p2[51:24]}};
        p_Val2_469_reg_42177 <= p_Val2_469_fu_21850_p2;
        p_Val2_471_reg_42010 <= {{r_V_100_fu_534_p2[44:24]}};
        p_Val2_472_reg_42192 <= p_Val2_472_fu_21979_p2;
        p_Val2_474_reg_42039 <= {{r_V_101_fu_478_p2[42:24]}};
        p_Val2_475_reg_42207 <= p_Val2_475_fu_22108_p2;
        p_Val2_477_reg_42068 <= {{r_V_102_fu_474_p2[40:24]}};
        p_Val2_478_reg_42222 <= p_Val2_478_fu_22237_p2;
        p_Val2_480_reg_42097 <= {{r_V_103_fu_469_p2[46:24]}};
        p_Val2_481_reg_42237 <= p_Val2_481_fu_22366_p2;
        p_Val2_484_reg_42264 <= p_Val2_484_fu_22548_p2;
        p_Val2_487_reg_42295 <= p_Val2_487_fu_22612_p2;
        p_Val2_490_reg_42326 <= p_Val2_490_fu_22676_p2;
        p_Val2_493_reg_42357 <= p_Val2_493_fu_22740_p2;
        p_Val2_496_reg_42388 <= p_Val2_496_fu_22804_p2;
        p_Val2_499_reg_42419 <= p_Val2_499_fu_22868_p2;
        p_Val2_502_reg_42438 <= p_Val2_502_fu_22951_p2;
        p_Val2_505_reg_42465 <= p_Val2_505_fu_23131_p2;
        p_Val2_508_reg_42496 <= p_Val2_508_fu_23195_p2;
        p_Val2_510_reg_42521 <= {{r_V_113_fu_535_p2[54:24]}};
        p_Val2_513_reg_42550 <= {{r_V_114_fu_475_p2[41:24]}};
        p_Val2_516_reg_42579 <= {{r_V_115_fu_468_p2[44:24]}};
        p_Val2_519_reg_42608 <= {{r_V_116_fu_537_p2[44:24]}};
        p_Val2_522_reg_42637 <= {{r_V_117_fu_519_p2[46:24]}};
        p_Val2_525_reg_42666 <= {{r_V_118_fu_470_p2[42:24]}};
        p_Val2_528_reg_42695 <= {{r_V_119_fu_542_p2[44:24]}};
        p_Val2_531_reg_42724 <= {{r_V_120_fu_520_p2[43:24]}};
        p_Val2_534_reg_42753 <= {{r_V_121_fu_477_p2[43:24]}};
        p_Val2_538_reg_42830 <= p_Val2_538_fu_27979_p2;
        p_Val2_541_reg_42857 <= p_Val2_541_fu_28159_p2;
        p_Val2_544_reg_42888 <= p_Val2_544_fu_28223_p2;
        p_Val2_547_reg_42919 <= p_Val2_547_fu_28287_p2;
        p_Val2_550_reg_42950 <= p_Val2_550_fu_28351_p2;
        p_Val2_553_reg_42981 <= p_Val2_553_fu_28415_p2;
        p_Val2_556_reg_43012 <= p_Val2_556_fu_28479_p2;
        p_Val2_559_reg_43043 <= p_Val2_559_fu_28543_p2;
        p_Val2_562_reg_43074 <= p_Val2_562_fu_28607_p2;
        p_Val2_564_reg_43099 <= {{r_V_131_fu_506_p2[43:24]}};
        p_Val2_567_reg_43128 <= {{r_V_132_fu_533_p2[42:24]}};
        p_Val2_570_reg_43157 <= {{r_V_133_fu_486_p2[42:24]}};
        p_Val2_573_reg_43186 <= {{r_V_134_fu_525_p2[43:24]}};
        p_Val2_576_reg_43215 <= {{r_V_135_fu_496_p2[42:24]}};
        p_Val2_579_reg_43244 <= {{r_V_136_fu_500_p2[42:24]}};
        p_Val2_582_reg_43273 <= {{r_V_137_fu_464_p2[40:24]}};
        p_Val2_585_reg_43302 <= {{r_V_138_fu_528_p2[41:24]}};
        p_Val2_589_reg_43325 <= p_Val2_589_fu_29046_p2;
        p_Val2_592_reg_43532 <= p_Val2_592_fu_33614_p2;
        p_Val2_595_reg_43563 <= p_Val2_595_fu_33678_p2;
        p_Val2_598_reg_43594 <= p_Val2_598_fu_33742_p2;
        p_Val2_601_reg_43625 <= p_Val2_601_fu_33806_p2;
        p_Val2_604_reg_43656 <= p_Val2_604_fu_33870_p2;
        p_Val2_607_reg_43687 <= p_Val2_607_fu_33934_p2;
        p_Val2_610_reg_43718 <= p_Val2_610_fu_33998_p2;
        p_Val2_613_reg_43749 <= p_Val2_613_fu_34062_p2;
        p_Val2_616_reg_43780 <= p_Val2_616_fu_34126_p2;
        p_Val2_618_reg_43805 <= {{r_V_149_fu_493_p2[54:24]}};
        p_Val2_621_reg_43834 <= {{r_V_150_fu_531_p2[41:24]}};
        p_Val2_624_reg_43863 <= {{r_V_151_fu_517_p2[43:24]}};
        p_Val2_627_reg_43892 <= {{r_V_152_fu_516_p2[49:24]}};
        p_Val2_630_reg_43921 <= {{r_V_153_fu_473_p2[49:24]}};
        p_Val2_633_reg_43950 <= {{r_V_154_fu_523_p2[41:24]}};
        p_Val2_636_reg_43979 <= {{r_V_155_fu_483_p2[43:24]}};
        p_Val2_640_reg_44002 <= p_Val2_640_fu_34538_p2;
        p_Val2_642_reg_44023 <= {{r_V_157_fu_467_p2[49:24]}};
        p_Val2_717_reg_43347 <= p_Val2_717_fu_31020_p2;
        p_Val2_719_reg_43367 <= p_Val2_719_fu_31056_p2;
        p_Val2_721_reg_43387 <= p_Val2_721_fu_31092_p2;
        p_Val2_723_reg_43407 <= p_Val2_723_fu_31128_p2;
        p_Val2_725_reg_43427 <= p_Val2_725_fu_31164_p2;
        p_Val2_727_reg_43447 <= p_Val2_727_fu_31200_p2;
        p_Val2_729_reg_43467 <= p_Val2_729_fu_31236_p2;
        p_Val2_731_reg_43487 <= p_Val2_731_fu_31272_p2;
        p_Val2_733_reg_43507 <= p_Val2_733_fu_31308_p2;
        p_read_27_reg_41274 <= p_read8_int_reg;
        p_read_27_reg_41274_pp0_iter1_reg <= p_read_27_reg_41274;
        p_read_27_reg_41274_pp0_iter2_reg <= p_read_27_reg_41274_pp0_iter1_reg;
        p_read_28_reg_41284 <= p_read7_int_reg;
        p_read_28_reg_41284_pp0_iter1_reg <= p_read_28_reg_41284;
        p_read_28_reg_41284_pp0_iter2_reg <= p_read_28_reg_41284_pp0_iter1_reg;
        p_read_29_reg_41293 <= p_read6_int_reg;
        p_read_29_reg_41293_pp0_iter1_reg <= p_read_29_reg_41293;
        p_read_30_reg_41303 <= p_read5_int_reg;
        p_read_30_reg_41303_pp0_iter1_reg <= p_read_30_reg_41303;
        p_read_31_reg_41314 <= p_read4_int_reg;
        p_read_32_reg_41324 <= p_read3_int_reg;
        r_V_100_reg_9159 <= r_V_100_fu_534_p2;
        r_V_101_reg_9163 <= r_V_101_fu_478_p2;
        r_V_102_reg_9167 <= r_V_102_fu_474_p2;
        r_V_103_reg_9171 <= r_V_103_fu_469_p2;
        r_V_104_reg_12983 <= r_V_104_fu_466_p2;
        r_V_105_reg_12987 <= r_V_105_fu_539_p2;
        r_V_106_reg_12991 <= r_V_106_fu_512_p2;
        r_V_107_reg_12995 <= r_V_107_fu_463_p2;
        r_V_108_reg_12999 <= r_V_108_fu_529_p2;
        r_V_109_reg_13003 <= r_V_109_fu_485_p2;
        r_V_111_reg_13007 <= r_V_111_fu_526_p2;
        r_V_112_reg_13011 <= r_V_112_fu_471_p2;
        r_V_113_reg_13015 <= r_V_113_fu_535_p2;
        r_V_114_reg_13019 <= r_V_114_fu_475_p2;
        r_V_115_reg_13023 <= r_V_115_fu_468_p2;
        r_V_116_reg_13027 <= r_V_116_fu_537_p2;
        r_V_117_reg_13031 <= r_V_117_fu_519_p2;
        r_V_118_reg_13035 <= r_V_118_fu_470_p2;
        r_V_119_reg_13039 <= r_V_119_fu_542_p2;
        r_V_120_reg_13043 <= r_V_120_fu_520_p2;
        r_V_121_reg_13047 <= r_V_121_fu_477_p2;
        r_V_123_reg_15547 <= r_V_123_fu_472_p2;
        r_V_124_reg_15551 <= r_V_124_fu_462_p2;
        r_V_125_reg_15555 <= r_V_125_fu_510_p2;
        r_V_126_reg_15559 <= r_V_126_fu_515_p2;
        r_V_127_reg_15563 <= r_V_127_fu_479_p2;
        r_V_128_reg_15567 <= r_V_128_fu_513_p2;
        r_V_129_reg_15571 <= r_V_129_fu_521_p2;
        r_V_130_reg_15575 <= r_V_130_fu_491_p2;
        r_V_131_reg_15579 <= r_V_131_fu_506_p2;
        r_V_132_reg_15583 <= r_V_132_fu_533_p2;
        r_V_133_reg_15587 <= r_V_133_fu_486_p2;
        r_V_134_reg_15591 <= r_V_134_fu_525_p2;
        r_V_135_reg_15595 <= r_V_135_fu_496_p2;
        r_V_136_reg_15599 <= r_V_136_fu_500_p2;
        r_V_137_reg_15603 <= r_V_137_fu_464_p2;
        r_V_138_reg_15607 <= r_V_138_fu_528_p2;
        r_V_140_reg_17175 <= r_V_140_fu_481_p2;
        r_V_141_reg_17179 <= r_V_141_fu_541_p2;
        r_V_142_reg_17183 <= r_V_142_fu_492_p2;
        r_V_143_reg_17187 <= r_V_143_fu_540_p2;
        r_V_144_reg_17191 <= r_V_144_fu_490_p2;
        r_V_145_reg_17195 <= r_V_145_fu_476_p2;
        r_V_146_reg_17199 <= r_V_146_fu_514_p2;
        r_V_147_reg_17203 <= r_V_147_fu_508_p2;
        r_V_148_reg_17207 <= r_V_148_fu_518_p2;
        r_V_149_reg_17211 <= r_V_149_fu_493_p2;
        r_V_150_reg_17215 <= r_V_150_fu_531_p2;
        r_V_151_reg_17219 <= r_V_151_fu_517_p2;
        r_V_152_reg_17223 <= r_V_152_fu_516_p2;
        r_V_153_reg_17227 <= r_V_153_fu_473_p2;
        r_V_154_reg_17231 <= r_V_154_fu_523_p2;
        r_V_155_reg_17235 <= r_V_155_fu_483_p2;
        r_V_157_reg_17239 <= r_V_157_fu_467_p2;
        r_V_78_reg_9075 <= r_V_78_fu_527_p2;
        r_V_79_reg_9079 <= r_V_79_fu_484_p2;
        r_V_80_reg_9083 <= r_V_80_fu_509_p2;
        r_V_81_reg_9087 <= r_V_81_fu_489_p2;
        r_V_82_reg_9091 <= r_V_82_fu_497_p2;
        r_V_83_reg_9095 <= r_V_83_fu_507_p2;
        r_V_84_reg_9099 <= r_V_84_fu_494_p2;
        r_V_85_reg_9103 <= r_V_85_fu_495_p2;
        r_V_86_reg_9107 <= r_V_86_fu_505_p2;
        r_V_87_reg_9111 <= r_V_87_fu_538_p2;
        r_V_88_reg_9115 <= r_V_88_fu_498_p2;
        r_V_89_reg_9119 <= r_V_89_fu_482_p2;
        r_V_90_reg_9123 <= r_V_90_fu_480_p2;
        r_V_92_reg_9127 <= r_V_92_fu_522_p2;
        r_V_93_reg_9131 <= r_V_93_fu_532_p2;
        r_V_94_reg_9135 <= r_V_94_fu_499_p2;
        r_V_95_reg_9139 <= r_V_95_fu_503_p2;
        r_V_96_reg_9143 <= r_V_96_fu_530_p2;
        r_V_97_reg_9147 <= r_V_97_fu_504_p2;
        r_V_98_reg_9151 <= r_V_98_fu_501_p2;
        r_V_99_reg_9155 <= r_V_99_fu_465_p2;
        r_V_reg_9071 <= r_V_fu_536_p2;
        rhs_101_reg_42171 <= rhs_101_fu_21836_p3;
        rhs_98_reg_42135 <= rhs_98_fu_21437_p3;
        tmp_1005_reg_43313 <= r_V_138_fu_528_p2[32'd23];
        tmp_1011_reg_42130 <= sub_ln823_3_fu_18952_p2[32'd23];
        tmp_1011_reg_42130_pp0_iter1_reg <= tmp_1011_reg_42130;
        tmp_1071_reg_43816 <= r_V_149_fu_493_p2[32'd23];
        tmp_1077_reg_43845 <= r_V_150_fu_531_p2[32'd23];
        tmp_1083_reg_43874 <= r_V_151_fu_517_p2[32'd23];
        tmp_1089_reg_43903 <= r_V_152_fu_516_p2[32'd23];
        tmp_1095_reg_43932 <= r_V_153_fu_473_p2[32'd23];
        tmp_1101_reg_43961 <= r_V_154_fu_523_p2[32'd23];
        tmp_1107_reg_43990 <= r_V_155_fu_483_p2[32'd23];
        tmp_1119_reg_44034 <= r_V_157_fu_467_p2[32'd23];
        tmp_693_reg_41629 <= r_V_86_fu_505_p2[32'd23];
        tmp_699_reg_41658 <= r_V_87_fu_538_p2[32'd23];
        tmp_705_reg_41687 <= r_V_88_fu_498_p2[32'd23];
        tmp_711_reg_41716 <= r_V_89_fu_482_p2[32'd23];
        tmp_717_reg_41745 <= r_V_90_fu_480_p2[32'd23];
        tmp_729_reg_41789 <= r_V_92_fu_522_p2[32'd23];
        tmp_735_reg_41818 <= r_V_93_fu_532_p2[32'd23];
        tmp_741_reg_41847 <= r_V_94_fu_499_p2[32'd23];
        tmp_747_reg_41876 <= r_V_95_fu_503_p2[32'd23];
        tmp_753_reg_41905 <= r_V_96_fu_530_p2[32'd23];
        tmp_759_reg_41934 <= r_V_97_fu_504_p2[32'd23];
        tmp_765_reg_41963 <= r_V_98_fu_501_p2[32'd23];
        tmp_771_reg_41992 <= r_V_99_fu_465_p2[32'd23];
        tmp_777_reg_42021 <= r_V_100_fu_534_p2[32'd23];
        tmp_783_reg_42050 <= r_V_101_fu_478_p2[32'd23];
        tmp_789_reg_42079 <= r_V_102_fu_474_p2[32'd23];
        tmp_795_reg_42108 <= r_V_103_fu_469_p2[32'd23];
        tmp_837_reg_42120 <= sub_ln823_fu_18876_p2[32'd23];
        tmp_855_reg_42532 <= r_V_113_fu_535_p2[32'd23];
        tmp_861_reg_42561 <= r_V_114_fu_475_p2[32'd23];
        tmp_867_reg_42590 <= r_V_115_fu_468_p2[32'd23];
        tmp_873_reg_42619 <= r_V_116_fu_537_p2[32'd23];
        tmp_879_reg_42648 <= r_V_117_fu_519_p2[32'd23];
        tmp_885_reg_42677 <= r_V_118_fu_470_p2[32'd23];
        tmp_891_reg_42706 <= r_V_119_fu_542_p2[32'd23];
        tmp_897_reg_42735 <= r_V_120_fu_520_p2[32'd23];
        tmp_903_reg_42764 <= r_V_121_fu_477_p2[32'd23];
        tmp_909_reg_42125 <= sub_ln823_2_fu_18914_p2[32'd23];
        tmp_909_reg_42125_pp0_iter1_reg <= tmp_909_reg_42125;
        tmp_963_reg_43110 <= r_V_131_fu_506_p2[32'd23];
        tmp_969_reg_43139 <= r_V_132_fu_533_p2[32'd23];
        tmp_975_reg_43168 <= r_V_133_fu_486_p2[32'd23];
        tmp_981_reg_43197 <= r_V_134_fu_525_p2[32'd23];
        tmp_987_reg_43226 <= r_V_135_fu_496_p2[32'd23];
        tmp_993_reg_43255 <= r_V_136_fu_500_p2[32'd23];
        tmp_999_reg_43284 <= r_V_137_fu_464_p2[32'd23];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= select_ln302_306_fu_40396_p3;
        ap_return_1_int_reg <= select_ln302_308_fu_40498_p3;
        ap_return_2_int_reg <= select_ln302_310_fu_40600_p3;
        ap_return_3_int_reg <= select_ln302_312_fu_40702_p3;
        ap_return_4_int_reg <= select_ln302_314_fu_40804_p3;
        ap_return_5_int_reg <= select_ln302_316_fu_40906_p3;
        ap_return_6_int_reg <= select_ln302_318_fu_41008_p3;
        ap_return_7_int_reg <= select_ln302_320_fu_41110_p3;
        ap_return_8_int_reg <= select_ln302_322_fu_41212_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        p_read1_int_reg <= p_read1;
        p_read2_int_reg <= p_read2;
        p_read3_int_reg <= p_read3;
        p_read4_int_reg <= p_read4;
        p_read5_int_reg <= p_read5;
        p_read6_int_reg <= p_read6;
        p_read7_int_reg <= p_read7;
        p_read8_int_reg <= p_read8;
        p_read_int_reg <= p_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = select_ln302_306_fu_40396_p3;
    end else begin
        ap_return_0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = select_ln302_308_fu_40498_p3;
    end else begin
        ap_return_1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = select_ln302_310_fu_40600_p3;
    end else begin
        ap_return_2 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = select_ln302_312_fu_40702_p3;
    end else begin
        ap_return_3 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = select_ln302_314_fu_40804_p3;
    end else begin
        ap_return_4 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = select_ln302_316_fu_40906_p3;
    end else begin
        ap_return_5 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = select_ln302_318_fu_41008_p3;
    end else begin
        ap_return_6 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = select_ln302_320_fu_41110_p3;
    end else begin
        ap_return_7 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = select_ln302_322_fu_41212_p3;
    end else begin
        ap_return_8 = 'bx;
    end
end

assign Range2_all_ones_111_fu_22977_p3 = r_V_110_fu_22912_p2[32'd38];

assign Range2_all_ones_123_fu_28005_p3 = r_V_122_fu_27940_p2[32'd40];

assign Range2_all_ones_140_fu_29072_p3 = r_V_139_fu_29007_p2[32'd40];

assign Range2_all_ones_157_fu_34564_p3 = r_V_156_fu_34490_p2[32'd35];

assign Range2_all_ones_92_fu_18195_p3 = r_V_91_fu_18121_p2[32'd39];

assign and_ln891_100_fu_21646_p2 = (carry_199_fu_21600_p2 & Range2_all_ones_98_reg_41939);

assign and_ln891_101_fu_21771_p2 = (carry_201_fu_21725_p2 & Range2_all_ones_99_reg_41968);

assign and_ln891_102_fu_21916_p2 = (carry_203_fu_21870_p2 & Range2_all_ones_100_reg_41997);

assign and_ln891_103_fu_22045_p2 = (carry_205_fu_21999_p2 & Range2_all_ones_101_reg_42026);

assign and_ln891_104_fu_22174_p2 = (carry_207_fu_22128_p2 & Range2_all_ones_102_reg_42055);

assign and_ln891_105_fu_22303_p2 = (carry_209_fu_22257_p2 & Range2_all_ones_103_reg_42084);

assign and_ln891_106_fu_22432_p2 = (carry_211_fu_22386_p2 & Range2_all_ones_104_reg_42113);

assign and_ln891_107_fu_25594_p2 = (carry_213_fu_25549_p2 & Range2_all_ones_105_reg_42276);

assign and_ln891_108_fu_25719_p2 = (carry_215_fu_25674_p2 & Range2_all_ones_106_reg_42307);

assign and_ln891_109_fu_25844_p2 = (carry_217_fu_25799_p2 & Range2_all_ones_107_reg_42338);

assign and_ln891_110_fu_25969_p2 = (carry_219_fu_25924_p2 & Range2_all_ones_108_reg_42369);

assign and_ln891_111_fu_26094_p2 = (carry_221_fu_26049_p2 & Range2_all_ones_109_reg_42400);

assign and_ln891_112_fu_26219_p2 = (carry_223_fu_26174_p2 & Range2_all_ones_110_reg_42431);

assign and_ln891_113_fu_23029_p2 = (carry_225_fu_22971_p2 & Range2_all_ones_111_fu_22977_p3);

assign and_ln891_114_fu_26361_p2 = (carry_227_fu_26316_p2 & Range2_all_ones_112_reg_42477);

assign and_ln891_115_fu_26486_p2 = (carry_229_fu_26441_p2 & Range2_all_ones_113_reg_42508);

assign and_ln891_116_fu_26630_p2 = (carry_231_fu_26584_p2 & Range2_all_ones_114_reg_42537);

assign and_ln891_117_fu_26779_p2 = (carry_233_fu_26733_p2 & Range2_all_ones_115_reg_42566);

assign and_ln891_118_fu_26928_p2 = (carry_235_fu_26882_p2 & Range2_all_ones_116_reg_42595);

assign and_ln891_119_fu_27077_p2 = (carry_237_fu_27031_p2 & Range2_all_ones_117_reg_42624);

assign and_ln891_120_fu_27226_p2 = (carry_239_fu_27180_p2 & Range2_all_ones_118_reg_42653);

assign and_ln891_121_fu_27375_p2 = (carry_241_fu_27329_p2 & Range2_all_ones_119_reg_42682);

assign and_ln891_122_fu_27524_p2 = (carry_243_fu_27478_p2 & Range2_all_ones_120_reg_42711);

assign and_ln891_123_fu_27673_p2 = (carry_245_fu_27627_p2 & Range2_all_ones_121_reg_42740);

assign and_ln891_124_fu_27822_p2 = (carry_247_fu_27776_p2 & Range2_all_ones_122_reg_42769);

assign and_ln891_125_fu_28057_p2 = (carry_249_fu_27999_p2 & Range2_all_ones_123_fu_28005_p3);

assign and_ln891_126_fu_31392_p2 = (carry_251_fu_31347_p2 & Range2_all_ones_124_reg_42869);

assign and_ln891_127_fu_31517_p2 = (carry_253_fu_31472_p2 & Range2_all_ones_125_reg_42900);

assign and_ln891_128_fu_31642_p2 = (carry_255_fu_31597_p2 & Range2_all_ones_126_reg_42931);

assign and_ln891_129_fu_31767_p2 = (carry_257_fu_31722_p2 & Range2_all_ones_127_reg_42962);

assign and_ln891_130_fu_31892_p2 = (carry_259_fu_31847_p2 & Range2_all_ones_128_reg_42993);

assign and_ln891_131_fu_32017_p2 = (carry_261_fu_31972_p2 & Range2_all_ones_129_reg_43024);

assign and_ln891_132_fu_32142_p2 = (carry_263_fu_32097_p2 & Range2_all_ones_130_reg_43055);

assign and_ln891_133_fu_32267_p2 = (carry_265_fu_32222_p2 & Range2_all_ones_131_reg_43086);

assign and_ln891_134_fu_32415_p2 = (carry_267_fu_32369_p2 & Range2_all_ones_132_reg_43115);

assign and_ln891_135_fu_32564_p2 = (carry_269_fu_32518_p2 & Range2_all_ones_133_reg_43144);

assign and_ln891_136_fu_32713_p2 = (carry_271_fu_32667_p2 & Range2_all_ones_134_reg_43173);

assign and_ln891_137_fu_32862_p2 = (carry_273_fu_32816_p2 & Range2_all_ones_135_reg_43202);

assign and_ln891_138_fu_33011_p2 = (carry_275_fu_32965_p2 & Range2_all_ones_136_reg_43231);

assign and_ln891_139_fu_33160_p2 = (carry_277_fu_33114_p2 & Range2_all_ones_137_reg_43260);

assign and_ln891_140_fu_33309_p2 = (carry_279_fu_33263_p2 & Range2_all_ones_138_reg_43289);

assign and_ln891_141_fu_33458_p2 = (carry_281_fu_33412_p2 & Range2_all_ones_139_reg_43318);

assign and_ln891_142_fu_29124_p2 = (carry_283_fu_29066_p2 & Range2_all_ones_140_fu_29072_p3);

assign and_ln891_143_fu_37126_p2 = (carry_285_fu_37081_p2 & Range2_all_ones_141_reg_43544);

assign and_ln891_144_fu_37250_p2 = (carry_287_fu_37205_p2 & Range2_all_ones_142_reg_43575);

assign and_ln891_145_fu_37375_p2 = (carry_289_fu_37330_p2 & Range2_all_ones_143_reg_43606);

assign and_ln891_146_fu_37500_p2 = (carry_291_fu_37455_p2 & Range2_all_ones_144_reg_43637);

assign and_ln891_147_fu_37625_p2 = (carry_293_fu_37580_p2 & Range2_all_ones_145_reg_43668);

assign and_ln891_148_fu_37750_p2 = (carry_295_fu_37705_p2 & Range2_all_ones_146_reg_43699);

assign and_ln891_149_fu_37875_p2 = (carry_297_fu_37830_p2 & Range2_all_ones_147_reg_43730);

assign and_ln891_150_fu_38000_p2 = (carry_299_fu_37955_p2 & Range2_all_ones_148_reg_43761);

assign and_ln891_151_fu_38125_p2 = (carry_301_fu_38080_p2 & Range2_all_ones_149_reg_43792);

assign and_ln891_152_fu_38269_p2 = (carry_303_fu_38223_p2 & Range2_all_ones_150_reg_43821);

assign and_ln891_153_fu_38418_p2 = (carry_305_fu_38372_p2 & Range2_all_ones_151_reg_43850);

assign and_ln891_154_fu_38567_p2 = (carry_307_fu_38521_p2 & Range2_all_ones_152_reg_43879);

assign and_ln891_155_fu_38716_p2 = (carry_309_fu_38670_p2 & Range2_all_ones_153_reg_43908);

assign and_ln891_156_fu_38865_p2 = (carry_311_fu_38819_p2 & Range2_all_ones_154_reg_43937);

assign and_ln891_157_fu_39014_p2 = (carry_313_fu_38968_p2 & Range2_all_ones_155_reg_43966);

assign and_ln891_158_fu_39163_p2 = (carry_315_fu_39117_p2 & Range2_all_ones_156_reg_43995);

assign and_ln891_159_fu_34616_p2 = (carry_317_fu_34558_p2 & Range2_all_ones_157_fu_34564_p3);

assign and_ln891_160_fu_39329_p2 = (carry_319_fu_39283_p2 & Range2_all_ones_158_reg_44039);

assign and_ln891_81_fu_19144_p2 = (carry_161_fu_19099_p2 & Range2_all_ones_79_reg_41388);

assign and_ln891_82_fu_19269_p2 = (carry_163_fu_19224_p2 & Range2_all_ones_80_reg_41419);

assign and_ln891_83_fu_19394_p2 = (carry_165_fu_19349_p2 & Range2_all_ones_81_reg_41450);

assign and_ln891_84_fu_19519_p2 = (carry_167_fu_19474_p2 & Range2_all_ones_82_reg_41481);

assign and_ln891_85_fu_19644_p2 = (carry_169_fu_19599_p2 & Range2_all_ones_83_reg_41512);

assign and_ln891_86_fu_19769_p2 = (carry_171_fu_19724_p2 & Range2_all_ones_84_reg_41543);

assign and_ln891_87_fu_19894_p2 = (carry_173_fu_19849_p2 & Range2_all_ones_85_reg_41574);

assign and_ln891_88_fu_20019_p2 = (carry_175_fu_19974_p2 & Range2_all_ones_86_reg_41605);

assign and_ln891_89_fu_20167_p2 = (carry_177_fu_20121_p2 & Range2_all_ones_87_reg_41634);

assign and_ln891_90_fu_20316_p2 = (carry_179_fu_20270_p2 & Range2_all_ones_88_reg_41663);

assign and_ln891_91_fu_20465_p2 = (carry_181_fu_20419_p2 & Range2_all_ones_89_reg_41692);

assign and_ln891_92_fu_20614_p2 = (carry_183_fu_20568_p2 & Range2_all_ones_90_reg_41721);

assign and_ln891_93_fu_20763_p2 = (carry_185_fu_20717_p2 & Range2_all_ones_91_reg_41750);

assign and_ln891_94_fu_18247_p2 = (carry_187_fu_18189_p2 & Range2_all_ones_92_fu_18195_p3);

assign and_ln891_95_fu_20929_p2 = (carry_189_fu_20883_p2 & Range2_all_ones_93_reg_41794);

assign and_ln891_96_fu_21078_p2 = (carry_191_fu_21032_p2 & Range2_all_ones_94_reg_41823);

assign and_ln891_97_fu_21227_p2 = (carry_193_fu_21181_p2 & Range2_all_ones_95_reg_41852);

assign and_ln891_98_fu_21372_p2 = (carry_195_fu_21326_p2 & Range2_all_ones_96_reg_41881);

assign and_ln891_99_fu_21517_p2 = (carry_197_fu_21471_p2 & Range2_all_ones_97_reg_41910);

assign and_ln891_fu_19019_p2 = (carry_159_fu_18974_p2 & Range2_all_ones_reg_41357);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign carry_159_fu_18974_p2 = (xor_ln896_fu_18969_p2 & p_Result_403_reg_41339);

assign carry_161_fu_19099_p2 = (xor_ln896_244_fu_19094_p2 & p_Result_406_reg_41370);

assign carry_163_fu_19224_p2 = (xor_ln896_246_fu_19219_p2 & p_Result_409_reg_41401);

assign carry_165_fu_19349_p2 = (xor_ln896_248_fu_19344_p2 & p_Result_412_reg_41432);

assign carry_167_fu_19474_p2 = (xor_ln896_250_fu_19469_p2 & p_Result_415_reg_41463);

assign carry_169_fu_19599_p2 = (xor_ln896_252_fu_19594_p2 & p_Result_418_reg_41494);

assign carry_171_fu_19724_p2 = (xor_ln896_254_fu_19719_p2 & p_Result_421_reg_41525);

assign carry_173_fu_19849_p2 = (xor_ln896_256_fu_19844_p2 & p_Result_424_reg_41556);

assign carry_175_fu_19974_p2 = (xor_ln896_258_fu_19969_p2 & p_Result_427_reg_41587);

assign carry_177_fu_20121_p2 = (xor_ln896_260_fu_20115_p2 & p_Result_430_reg_41623);

assign carry_179_fu_20270_p2 = (xor_ln896_262_fu_20264_p2 & p_Result_433_reg_41652);

assign carry_181_fu_20419_p2 = (xor_ln896_264_fu_20413_p2 & p_Result_436_reg_41681);

assign carry_183_fu_20568_p2 = (xor_ln896_266_fu_20562_p2 & p_Result_439_reg_41710);

assign carry_185_fu_20717_p2 = (xor_ln896_268_fu_20711_p2 & p_Result_442_reg_41739);

assign carry_187_fu_18189_p2 = (xor_ln896_270_fu_18183_p2 & p_Result_445_fu_18149_p3);

assign carry_189_fu_20883_p2 = (xor_ln896_272_fu_20877_p2 & p_Result_448_reg_41783);

assign carry_191_fu_21032_p2 = (xor_ln896_274_fu_21026_p2 & p_Result_451_reg_41812);

assign carry_193_fu_21181_p2 = (xor_ln896_276_fu_21175_p2 & p_Result_454_reg_41841);

assign carry_195_fu_21326_p2 = (xor_ln896_278_fu_21320_p2 & p_Result_457_reg_41870);

assign carry_197_fu_21471_p2 = (xor_ln896_280_fu_21465_p2 & p_Result_460_reg_41899);

assign carry_199_fu_21600_p2 = (xor_ln896_282_fu_21594_p2 & p_Result_463_reg_41928);

assign carry_201_fu_21725_p2 = (xor_ln896_284_fu_21719_p2 & p_Result_466_reg_41957);

assign carry_203_fu_21870_p2 = (xor_ln896_286_fu_21864_p2 & p_Result_469_reg_41986);

assign carry_205_fu_21999_p2 = (xor_ln896_288_fu_21993_p2 & p_Result_472_reg_42015);

assign carry_207_fu_22128_p2 = (xor_ln896_290_fu_22122_p2 & p_Result_475_reg_42044);

assign carry_209_fu_22257_p2 = (xor_ln896_292_fu_22251_p2 & p_Result_478_reg_42073);

assign carry_211_fu_22386_p2 = (xor_ln896_294_fu_22380_p2 & p_Result_481_reg_42102);

assign carry_213_fu_25549_p2 = (xor_ln896_296_fu_25544_p2 & p_Result_484_reg_42258);

assign carry_215_fu_25674_p2 = (xor_ln896_298_fu_25669_p2 & p_Result_487_reg_42289);

assign carry_217_fu_25799_p2 = (xor_ln896_300_fu_25794_p2 & p_Result_490_reg_42320);

assign carry_219_fu_25924_p2 = (xor_ln896_302_fu_25919_p2 & p_Result_493_reg_42351);

assign carry_221_fu_26049_p2 = (xor_ln896_304_fu_26044_p2 & p_Result_496_reg_42382);

assign carry_223_fu_26174_p2 = (xor_ln896_306_fu_26169_p2 & p_Result_499_reg_42413);

assign carry_225_fu_22971_p2 = (xor_ln896_308_fu_22965_p2 & p_Result_502_fu_22940_p3);

assign carry_227_fu_26316_p2 = (xor_ln896_310_fu_26311_p2 & p_Result_505_reg_42459);

assign carry_229_fu_26441_p2 = (xor_ln896_312_fu_26436_p2 & p_Result_508_reg_42490);

assign carry_231_fu_26584_p2 = (xor_ln896_314_fu_26578_p2 & p_Result_511_reg_42526);

assign carry_233_fu_26733_p2 = (xor_ln896_316_fu_26727_p2 & p_Result_514_reg_42555);

assign carry_235_fu_26882_p2 = (xor_ln896_318_fu_26876_p2 & p_Result_517_reg_42584);

assign carry_237_fu_27031_p2 = (xor_ln896_320_fu_27025_p2 & p_Result_520_reg_42613);

assign carry_239_fu_27180_p2 = (xor_ln896_322_fu_27174_p2 & p_Result_523_reg_42642);

assign carry_241_fu_27329_p2 = (xor_ln896_324_fu_27323_p2 & p_Result_526_reg_42671);

assign carry_243_fu_27478_p2 = (xor_ln896_326_fu_27472_p2 & p_Result_529_reg_42700);

assign carry_245_fu_27627_p2 = (xor_ln896_328_fu_27621_p2 & p_Result_532_reg_42729);

assign carry_247_fu_27776_p2 = (xor_ln896_330_fu_27770_p2 & p_Result_535_reg_42758);

assign carry_249_fu_27999_p2 = (xor_ln896_332_fu_27993_p2 & p_Result_538_fu_27968_p3);

assign carry_251_fu_31347_p2 = (xor_ln896_334_fu_31342_p2 & p_Result_541_reg_42851);

assign carry_253_fu_31472_p2 = (xor_ln896_336_fu_31467_p2 & p_Result_544_reg_42882);

assign carry_255_fu_31597_p2 = (xor_ln896_338_fu_31592_p2 & p_Result_547_reg_42913);

assign carry_257_fu_31722_p2 = (xor_ln896_340_fu_31717_p2 & p_Result_550_reg_42944);

assign carry_259_fu_31847_p2 = (xor_ln896_342_fu_31842_p2 & p_Result_553_reg_42975);

assign carry_261_fu_31972_p2 = (xor_ln896_344_fu_31967_p2 & p_Result_556_reg_43006);

assign carry_263_fu_32097_p2 = (xor_ln896_346_fu_32092_p2 & p_Result_559_reg_43037);

assign carry_265_fu_32222_p2 = (xor_ln896_348_fu_32217_p2 & p_Result_562_reg_43068);

assign carry_267_fu_32369_p2 = (xor_ln896_350_fu_32363_p2 & p_Result_565_reg_43104);

assign carry_269_fu_32518_p2 = (xor_ln896_352_fu_32512_p2 & p_Result_568_reg_43133);

assign carry_271_fu_32667_p2 = (xor_ln896_354_fu_32661_p2 & p_Result_571_reg_43162);

assign carry_273_fu_32816_p2 = (xor_ln896_356_fu_32810_p2 & p_Result_574_reg_43191);

assign carry_275_fu_32965_p2 = (xor_ln896_358_fu_32959_p2 & p_Result_577_reg_43220);

assign carry_277_fu_33114_p2 = (xor_ln896_360_fu_33108_p2 & p_Result_580_reg_43249);

assign carry_279_fu_33263_p2 = (xor_ln896_362_fu_33257_p2 & p_Result_583_reg_43278);

assign carry_281_fu_33412_p2 = (xor_ln896_364_fu_33406_p2 & p_Result_586_reg_43307);

assign carry_283_fu_29066_p2 = (xor_ln896_366_fu_29060_p2 & p_Result_589_fu_29035_p3);

assign carry_285_fu_37081_p2 = (xor_ln896_368_fu_37076_p2 & p_Result_592_reg_43526);

assign carry_287_fu_37205_p2 = (xor_ln896_370_fu_37200_p2 & p_Result_595_reg_43557);

assign carry_289_fu_37330_p2 = (xor_ln896_372_fu_37325_p2 & p_Result_598_reg_43588);

assign carry_291_fu_37455_p2 = (xor_ln896_374_fu_37450_p2 & p_Result_601_reg_43619);

assign carry_293_fu_37580_p2 = (xor_ln896_376_fu_37575_p2 & p_Result_604_reg_43650);

assign carry_295_fu_37705_p2 = (xor_ln896_378_fu_37700_p2 & p_Result_607_reg_43681);

assign carry_297_fu_37830_p2 = (xor_ln896_380_fu_37825_p2 & p_Result_610_reg_43712);

assign carry_299_fu_37955_p2 = (xor_ln896_382_fu_37950_p2 & p_Result_613_reg_43743);

assign carry_301_fu_38080_p2 = (xor_ln896_384_fu_38075_p2 & p_Result_616_reg_43774);

assign carry_303_fu_38223_p2 = (xor_ln896_386_fu_38217_p2 & p_Result_619_reg_43810);

assign carry_305_fu_38372_p2 = (xor_ln896_388_fu_38366_p2 & p_Result_622_reg_43839);

assign carry_307_fu_38521_p2 = (xor_ln896_390_fu_38515_p2 & p_Result_625_reg_43868);

assign carry_309_fu_38670_p2 = (xor_ln896_392_fu_38664_p2 & p_Result_628_reg_43897);

assign carry_311_fu_38819_p2 = (xor_ln896_394_fu_38813_p2 & p_Result_631_reg_43926);

assign carry_313_fu_38968_p2 = (xor_ln896_396_fu_38962_p2 & p_Result_634_reg_43955);

assign carry_315_fu_39117_p2 = (xor_ln896_398_fu_39111_p2 & p_Result_637_reg_43984);

assign carry_317_fu_34558_p2 = (xor_ln896_400_fu_34552_p2 & p_Result_640_fu_34518_p3);

assign carry_319_fu_39283_p2 = (xor_ln896_402_fu_39277_p2 & p_Result_643_reg_44028);

assign deleted_ones_162_fu_19139_p2 = (or_ln890_81_fu_19133_p2 & Range2_all_ones_79_reg_41388);

assign deleted_ones_163_fu_19264_p2 = (or_ln890_82_fu_19258_p2 & Range2_all_ones_80_reg_41419);

assign deleted_ones_164_fu_19389_p2 = (or_ln890_83_fu_19383_p2 & Range2_all_ones_81_reg_41450);

assign deleted_ones_165_fu_19514_p2 = (or_ln890_84_fu_19508_p2 & Range2_all_ones_82_reg_41481);

assign deleted_ones_166_fu_19639_p2 = (or_ln890_85_fu_19633_p2 & Range2_all_ones_83_reg_41512);

assign deleted_ones_167_fu_19764_p2 = (or_ln890_86_fu_19758_p2 & Range2_all_ones_84_reg_41543);

assign deleted_ones_168_fu_19889_p2 = (or_ln890_87_fu_19883_p2 & Range2_all_ones_85_reg_41574);

assign deleted_ones_169_fu_20014_p2 = (or_ln890_88_fu_20008_p2 & Range2_all_ones_86_reg_41605);

assign deleted_ones_170_fu_20162_p2 = (or_ln890_89_fu_20156_p2 & Range2_all_ones_87_reg_41634);

assign deleted_ones_171_fu_20311_p2 = (or_ln890_90_fu_20305_p2 & Range2_all_ones_88_reg_41663);

assign deleted_ones_172_fu_20460_p2 = (or_ln890_91_fu_20454_p2 & Range2_all_ones_89_reg_41692);

assign deleted_ones_173_fu_20609_p2 = (or_ln890_92_fu_20603_p2 & Range2_all_ones_90_reg_41721);

assign deleted_ones_174_fu_20758_p2 = (or_ln890_93_fu_20752_p2 & Range2_all_ones_91_reg_41750);

assign deleted_ones_175_fu_18241_p2 = (or_ln890_94_fu_18235_p2 & Range2_all_ones_92_fu_18195_p3);

assign deleted_ones_176_fu_20924_p2 = (or_ln890_95_fu_20918_p2 & Range2_all_ones_93_reg_41794);

assign deleted_ones_177_fu_21073_p2 = (or_ln890_96_fu_21067_p2 & Range2_all_ones_94_reg_41823);

assign deleted_ones_178_fu_21222_p2 = (or_ln890_97_fu_21216_p2 & Range2_all_ones_95_reg_41852);

assign deleted_ones_179_fu_21367_p2 = (or_ln890_98_fu_21361_p2 & Range2_all_ones_96_reg_41881);

assign deleted_ones_180_fu_21512_p2 = (or_ln890_99_fu_21506_p2 & Range2_all_ones_97_reg_41910);

assign deleted_ones_181_fu_21641_p2 = (or_ln890_100_fu_21635_p2 & Range2_all_ones_98_reg_41939);

assign deleted_ones_182_fu_21766_p2 = (or_ln890_101_fu_21760_p2 & Range2_all_ones_99_reg_41968);

assign deleted_ones_183_fu_21911_p2 = (or_ln890_102_fu_21905_p2 & Range2_all_ones_100_reg_41997);

assign deleted_ones_184_fu_22040_p2 = (or_ln890_103_fu_22034_p2 & Range2_all_ones_101_reg_42026);

assign deleted_ones_185_fu_22169_p2 = (or_ln890_104_fu_22163_p2 & Range2_all_ones_102_reg_42055);

assign deleted_ones_186_fu_22298_p2 = (or_ln890_105_fu_22292_p2 & Range2_all_ones_103_reg_42084);

assign deleted_ones_187_fu_22427_p2 = (or_ln890_106_fu_22421_p2 & Range2_all_ones_104_reg_42113);

assign deleted_ones_188_fu_25589_p2 = (or_ln890_107_fu_25583_p2 & Range2_all_ones_105_reg_42276);

assign deleted_ones_189_fu_25714_p2 = (or_ln890_108_fu_25708_p2 & Range2_all_ones_106_reg_42307);

assign deleted_ones_190_fu_25839_p2 = (or_ln890_109_fu_25833_p2 & Range2_all_ones_107_reg_42338);

assign deleted_ones_191_fu_25964_p2 = (or_ln890_110_fu_25958_p2 & Range2_all_ones_108_reg_42369);

assign deleted_ones_192_fu_26089_p2 = (or_ln890_111_fu_26083_p2 & Range2_all_ones_109_reg_42400);

assign deleted_ones_193_fu_26214_p2 = (or_ln890_112_fu_26208_p2 & Range2_all_ones_110_reg_42431);

assign deleted_ones_194_fu_23023_p2 = (or_ln890_113_fu_23017_p2 & Range2_all_ones_111_fu_22977_p3);

assign deleted_ones_195_fu_26356_p2 = (or_ln890_114_fu_26350_p2 & Range2_all_ones_112_reg_42477);

assign deleted_ones_196_fu_26481_p2 = (or_ln890_115_fu_26475_p2 & Range2_all_ones_113_reg_42508);

assign deleted_ones_197_fu_26625_p2 = (or_ln890_116_fu_26619_p2 & Range2_all_ones_114_reg_42537);

assign deleted_ones_198_fu_26774_p2 = (or_ln890_117_fu_26768_p2 & Range2_all_ones_115_reg_42566);

assign deleted_ones_199_fu_26923_p2 = (or_ln890_118_fu_26917_p2 & Range2_all_ones_116_reg_42595);

assign deleted_ones_200_fu_27072_p2 = (or_ln890_119_fu_27066_p2 & Range2_all_ones_117_reg_42624);

assign deleted_ones_201_fu_27221_p2 = (or_ln890_120_fu_27215_p2 & Range2_all_ones_118_reg_42653);

assign deleted_ones_202_fu_27370_p2 = (or_ln890_121_fu_27364_p2 & Range2_all_ones_119_reg_42682);

assign deleted_ones_203_fu_27519_p2 = (or_ln890_122_fu_27513_p2 & Range2_all_ones_120_reg_42711);

assign deleted_ones_204_fu_27668_p2 = (or_ln890_123_fu_27662_p2 & Range2_all_ones_121_reg_42740);

assign deleted_ones_205_fu_27817_p2 = (or_ln890_124_fu_27811_p2 & Range2_all_ones_122_reg_42769);

assign deleted_ones_206_fu_28051_p2 = (or_ln890_125_fu_28045_p2 & Range2_all_ones_123_fu_28005_p3);

assign deleted_ones_207_fu_31387_p2 = (or_ln890_126_fu_31381_p2 & Range2_all_ones_124_reg_42869);

assign deleted_ones_208_fu_31512_p2 = (or_ln890_127_fu_31506_p2 & Range2_all_ones_125_reg_42900);

assign deleted_ones_209_fu_31637_p2 = (or_ln890_128_fu_31631_p2 & Range2_all_ones_126_reg_42931);

assign deleted_ones_210_fu_31762_p2 = (or_ln890_129_fu_31756_p2 & Range2_all_ones_127_reg_42962);

assign deleted_ones_211_fu_31887_p2 = (or_ln890_130_fu_31881_p2 & Range2_all_ones_128_reg_42993);

assign deleted_ones_212_fu_32012_p2 = (or_ln890_131_fu_32006_p2 & Range2_all_ones_129_reg_43024);

assign deleted_ones_213_fu_32137_p2 = (or_ln890_132_fu_32131_p2 & Range2_all_ones_130_reg_43055);

assign deleted_ones_214_fu_32262_p2 = (or_ln890_133_fu_32256_p2 & Range2_all_ones_131_reg_43086);

assign deleted_ones_215_fu_32410_p2 = (or_ln890_134_fu_32404_p2 & Range2_all_ones_132_reg_43115);

assign deleted_ones_216_fu_32559_p2 = (or_ln890_135_fu_32553_p2 & Range2_all_ones_133_reg_43144);

assign deleted_ones_217_fu_32708_p2 = (or_ln890_136_fu_32702_p2 & Range2_all_ones_134_reg_43173);

assign deleted_ones_218_fu_32857_p2 = (or_ln890_137_fu_32851_p2 & Range2_all_ones_135_reg_43202);

assign deleted_ones_219_fu_33006_p2 = (or_ln890_138_fu_33000_p2 & Range2_all_ones_136_reg_43231);

assign deleted_ones_220_fu_33155_p2 = (or_ln890_139_fu_33149_p2 & Range2_all_ones_137_reg_43260);

assign deleted_ones_221_fu_33304_p2 = (or_ln890_140_fu_33298_p2 & Range2_all_ones_138_reg_43289);

assign deleted_ones_222_fu_33453_p2 = (or_ln890_141_fu_33447_p2 & Range2_all_ones_139_reg_43318);

assign deleted_ones_223_fu_29118_p2 = (or_ln890_142_fu_29112_p2 & Range2_all_ones_140_fu_29072_p3);

assign deleted_ones_224_fu_37121_p2 = (or_ln890_143_fu_37115_p2 & Range2_all_ones_141_reg_43544);

assign deleted_ones_225_fu_37245_p2 = (or_ln890_144_fu_37239_p2 & Range2_all_ones_142_reg_43575);

assign deleted_ones_226_fu_37370_p2 = (or_ln890_145_fu_37364_p2 & Range2_all_ones_143_reg_43606);

assign deleted_ones_227_fu_37495_p2 = (or_ln890_146_fu_37489_p2 & Range2_all_ones_144_reg_43637);

assign deleted_ones_228_fu_37620_p2 = (or_ln890_147_fu_37614_p2 & Range2_all_ones_145_reg_43668);

assign deleted_ones_229_fu_37745_p2 = (or_ln890_148_fu_37739_p2 & Range2_all_ones_146_reg_43699);

assign deleted_ones_230_fu_37870_p2 = (or_ln890_149_fu_37864_p2 & Range2_all_ones_147_reg_43730);

assign deleted_ones_231_fu_37995_p2 = (or_ln890_150_fu_37989_p2 & Range2_all_ones_148_reg_43761);

assign deleted_ones_232_fu_38120_p2 = (or_ln890_151_fu_38114_p2 & Range2_all_ones_149_reg_43792);

assign deleted_ones_233_fu_38264_p2 = (or_ln890_152_fu_38258_p2 & Range2_all_ones_150_reg_43821);

assign deleted_ones_234_fu_38413_p2 = (or_ln890_153_fu_38407_p2 & Range2_all_ones_151_reg_43850);

assign deleted_ones_235_fu_38562_p2 = (or_ln890_154_fu_38556_p2 & Range2_all_ones_152_reg_43879);

assign deleted_ones_236_fu_38711_p2 = (or_ln890_155_fu_38705_p2 & Range2_all_ones_153_reg_43908);

assign deleted_ones_237_fu_38860_p2 = (or_ln890_156_fu_38854_p2 & Range2_all_ones_154_reg_43937);

assign deleted_ones_238_fu_39009_p2 = (or_ln890_157_fu_39003_p2 & Range2_all_ones_155_reg_43966);

assign deleted_ones_239_fu_39158_p2 = (or_ln890_158_fu_39152_p2 & Range2_all_ones_156_reg_43995);

assign deleted_ones_240_fu_34610_p2 = (or_ln890_159_fu_34604_p2 & Range2_all_ones_157_fu_34564_p3);

assign deleted_ones_241_fu_39324_p2 = (or_ln890_160_fu_39318_p2 & Range2_all_ones_158_reg_44039);

assign deleted_ones_fu_19014_p2 = (or_ln890_fu_19008_p2 & Range2_all_ones_reg_41357);

assign deleted_zeros_100_fu_22015_p2 = (or_ln888_103_fu_22009_p2 ^ Range2_all_ones_101_reg_42026);

assign deleted_zeros_101_fu_22144_p2 = (or_ln888_104_fu_22138_p2 ^ Range2_all_ones_102_reg_42055);

assign deleted_zeros_102_fu_22273_p2 = (or_ln888_105_fu_22267_p2 ^ Range2_all_ones_103_reg_42084);

assign deleted_zeros_103_fu_22402_p2 = (or_ln888_106_fu_22396_p2 ^ Range2_all_ones_104_reg_42113);

assign deleted_zeros_104_fu_25564_p2 = (or_ln888_107_fu_25559_p2 ^ Range2_all_ones_105_reg_42276);

assign deleted_zeros_105_fu_25689_p2 = (or_ln888_108_fu_25684_p2 ^ Range2_all_ones_106_reg_42307);

assign deleted_zeros_106_fu_25814_p2 = (or_ln888_109_fu_25809_p2 ^ Range2_all_ones_107_reg_42338);

assign deleted_zeros_107_fu_25939_p2 = (or_ln888_110_fu_25934_p2 ^ Range2_all_ones_108_reg_42369);

assign deleted_zeros_108_fu_26064_p2 = (or_ln888_111_fu_26059_p2 ^ Range2_all_ones_109_reg_42400);

assign deleted_zeros_109_fu_26189_p2 = (or_ln888_112_fu_26184_p2 ^ Range2_all_ones_110_reg_42431);

assign deleted_zeros_110_fu_22997_p2 = (or_ln888_113_fu_22991_p2 ^ Range2_all_ones_111_fu_22977_p3);

assign deleted_zeros_111_fu_26331_p2 = (or_ln888_114_fu_26326_p2 ^ Range2_all_ones_112_reg_42477);

assign deleted_zeros_112_fu_26456_p2 = (or_ln888_115_fu_26451_p2 ^ Range2_all_ones_113_reg_42508);

assign deleted_zeros_113_fu_26600_p2 = (or_ln888_116_fu_26594_p2 ^ Range2_all_ones_114_reg_42537);

assign deleted_zeros_114_fu_26749_p2 = (or_ln888_117_fu_26743_p2 ^ Range2_all_ones_115_reg_42566);

assign deleted_zeros_115_fu_26898_p2 = (or_ln888_118_fu_26892_p2 ^ Range2_all_ones_116_reg_42595);

assign deleted_zeros_116_fu_27047_p2 = (or_ln888_119_fu_27041_p2 ^ Range2_all_ones_117_reg_42624);

assign deleted_zeros_117_fu_27196_p2 = (or_ln888_120_fu_27190_p2 ^ Range2_all_ones_118_reg_42653);

assign deleted_zeros_118_fu_27345_p2 = (or_ln888_121_fu_27339_p2 ^ Range2_all_ones_119_reg_42682);

assign deleted_zeros_119_fu_27494_p2 = (or_ln888_122_fu_27488_p2 ^ Range2_all_ones_120_reg_42711);

assign deleted_zeros_120_fu_27643_p2 = (or_ln888_123_fu_27637_p2 ^ Range2_all_ones_121_reg_42740);

assign deleted_zeros_121_fu_27792_p2 = (or_ln888_124_fu_27786_p2 ^ Range2_all_ones_122_reg_42769);

assign deleted_zeros_122_fu_28025_p2 = (or_ln888_125_fu_28019_p2 ^ Range2_all_ones_123_fu_28005_p3);

assign deleted_zeros_123_fu_31362_p2 = (or_ln888_126_fu_31357_p2 ^ Range2_all_ones_124_reg_42869);

assign deleted_zeros_124_fu_31487_p2 = (or_ln888_127_fu_31482_p2 ^ Range2_all_ones_125_reg_42900);

assign deleted_zeros_125_fu_31612_p2 = (or_ln888_128_fu_31607_p2 ^ Range2_all_ones_126_reg_42931);

assign deleted_zeros_126_fu_31737_p2 = (or_ln888_129_fu_31732_p2 ^ Range2_all_ones_127_reg_42962);

assign deleted_zeros_127_fu_31862_p2 = (or_ln888_130_fu_31857_p2 ^ Range2_all_ones_128_reg_42993);

assign deleted_zeros_128_fu_31987_p2 = (or_ln888_131_fu_31982_p2 ^ Range2_all_ones_129_reg_43024);

assign deleted_zeros_129_fu_32112_p2 = (or_ln888_132_fu_32107_p2 ^ Range2_all_ones_130_reg_43055);

assign deleted_zeros_130_fu_32237_p2 = (or_ln888_133_fu_32232_p2 ^ Range2_all_ones_131_reg_43086);

assign deleted_zeros_131_fu_32385_p2 = (or_ln888_134_fu_32379_p2 ^ Range2_all_ones_132_reg_43115);

assign deleted_zeros_132_fu_32534_p2 = (or_ln888_135_fu_32528_p2 ^ Range2_all_ones_133_reg_43144);

assign deleted_zeros_133_fu_32683_p2 = (or_ln888_136_fu_32677_p2 ^ Range2_all_ones_134_reg_43173);

assign deleted_zeros_134_fu_32832_p2 = (or_ln888_137_fu_32826_p2 ^ Range2_all_ones_135_reg_43202);

assign deleted_zeros_135_fu_32981_p2 = (or_ln888_138_fu_32975_p2 ^ Range2_all_ones_136_reg_43231);

assign deleted_zeros_136_fu_33130_p2 = (or_ln888_139_fu_33124_p2 ^ Range2_all_ones_137_reg_43260);

assign deleted_zeros_137_fu_33279_p2 = (or_ln888_140_fu_33273_p2 ^ Range2_all_ones_138_reg_43289);

assign deleted_zeros_138_fu_33428_p2 = (or_ln888_141_fu_33422_p2 ^ Range2_all_ones_139_reg_43318);

assign deleted_zeros_139_fu_29092_p2 = (or_ln888_142_fu_29086_p2 ^ Range2_all_ones_140_fu_29072_p3);

assign deleted_zeros_140_fu_37096_p2 = (or_ln888_143_fu_37091_p2 ^ Range2_all_ones_141_reg_43544);

assign deleted_zeros_141_fu_37220_p2 = (or_ln888_144_fu_37215_p2 ^ Range2_all_ones_142_reg_43575);

assign deleted_zeros_142_fu_37345_p2 = (or_ln888_145_fu_37340_p2 ^ Range2_all_ones_143_reg_43606);

assign deleted_zeros_143_fu_37470_p2 = (or_ln888_146_fu_37465_p2 ^ Range2_all_ones_144_reg_43637);

assign deleted_zeros_144_fu_37595_p2 = (or_ln888_147_fu_37590_p2 ^ Range2_all_ones_145_reg_43668);

assign deleted_zeros_145_fu_37720_p2 = (or_ln888_148_fu_37715_p2 ^ Range2_all_ones_146_reg_43699);

assign deleted_zeros_146_fu_37845_p2 = (or_ln888_149_fu_37840_p2 ^ Range2_all_ones_147_reg_43730);

assign deleted_zeros_147_fu_37970_p2 = (or_ln888_150_fu_37965_p2 ^ Range2_all_ones_148_reg_43761);

assign deleted_zeros_148_fu_38095_p2 = (or_ln888_151_fu_38090_p2 ^ Range2_all_ones_149_reg_43792);

assign deleted_zeros_149_fu_38239_p2 = (or_ln888_152_fu_38233_p2 ^ Range2_all_ones_150_reg_43821);

assign deleted_zeros_150_fu_38388_p2 = (or_ln888_153_fu_38382_p2 ^ Range2_all_ones_151_reg_43850);

assign deleted_zeros_151_fu_38537_p2 = (or_ln888_154_fu_38531_p2 ^ Range2_all_ones_152_reg_43879);

assign deleted_zeros_152_fu_38686_p2 = (or_ln888_155_fu_38680_p2 ^ Range2_all_ones_153_reg_43908);

assign deleted_zeros_153_fu_38835_p2 = (or_ln888_156_fu_38829_p2 ^ Range2_all_ones_154_reg_43937);

assign deleted_zeros_154_fu_38984_p2 = (or_ln888_157_fu_38978_p2 ^ Range2_all_ones_155_reg_43966);

assign deleted_zeros_155_fu_39133_p2 = (or_ln888_158_fu_39127_p2 ^ Range2_all_ones_156_reg_43995);

assign deleted_zeros_156_fu_34584_p2 = (or_ln888_159_fu_34578_p2 ^ Range2_all_ones_157_fu_34564_p3);

assign deleted_zeros_157_fu_39299_p2 = (or_ln888_160_fu_39293_p2 ^ Range2_all_ones_158_reg_44039);

assign deleted_zeros_78_fu_19114_p2 = (or_ln888_81_fu_19109_p2 ^ Range2_all_ones_79_reg_41388);

assign deleted_zeros_79_fu_19239_p2 = (or_ln888_82_fu_19234_p2 ^ Range2_all_ones_80_reg_41419);

assign deleted_zeros_80_fu_19364_p2 = (or_ln888_83_fu_19359_p2 ^ Range2_all_ones_81_reg_41450);

assign deleted_zeros_81_fu_19489_p2 = (or_ln888_84_fu_19484_p2 ^ Range2_all_ones_82_reg_41481);

assign deleted_zeros_82_fu_19614_p2 = (or_ln888_85_fu_19609_p2 ^ Range2_all_ones_83_reg_41512);

assign deleted_zeros_83_fu_19739_p2 = (or_ln888_86_fu_19734_p2 ^ Range2_all_ones_84_reg_41543);

assign deleted_zeros_84_fu_19864_p2 = (or_ln888_87_fu_19859_p2 ^ Range2_all_ones_85_reg_41574);

assign deleted_zeros_85_fu_19989_p2 = (or_ln888_88_fu_19984_p2 ^ Range2_all_ones_86_reg_41605);

assign deleted_zeros_86_fu_20137_p2 = (or_ln888_89_fu_20131_p2 ^ Range2_all_ones_87_reg_41634);

assign deleted_zeros_87_fu_20286_p2 = (or_ln888_90_fu_20280_p2 ^ Range2_all_ones_88_reg_41663);

assign deleted_zeros_88_fu_20435_p2 = (or_ln888_91_fu_20429_p2 ^ Range2_all_ones_89_reg_41692);

assign deleted_zeros_89_fu_20584_p2 = (or_ln888_92_fu_20578_p2 ^ Range2_all_ones_90_reg_41721);

assign deleted_zeros_90_fu_20733_p2 = (or_ln888_93_fu_20727_p2 ^ Range2_all_ones_91_reg_41750);

assign deleted_zeros_91_fu_18215_p2 = (or_ln888_94_fu_18209_p2 ^ Range2_all_ones_92_fu_18195_p3);

assign deleted_zeros_92_fu_20899_p2 = (or_ln888_95_fu_20893_p2 ^ Range2_all_ones_93_reg_41794);

assign deleted_zeros_93_fu_21048_p2 = (or_ln888_96_fu_21042_p2 ^ Range2_all_ones_94_reg_41823);

assign deleted_zeros_94_fu_21197_p2 = (or_ln888_97_fu_21191_p2 ^ Range2_all_ones_95_reg_41852);

assign deleted_zeros_95_fu_21342_p2 = (or_ln888_98_fu_21336_p2 ^ Range2_all_ones_96_reg_41881);

assign deleted_zeros_96_fu_21487_p2 = (or_ln888_99_fu_21481_p2 ^ Range2_all_ones_97_reg_41910);

assign deleted_zeros_97_fu_21616_p2 = (or_ln888_100_fu_21610_p2 ^ Range2_all_ones_98_reg_41939);

assign deleted_zeros_98_fu_21741_p2 = (or_ln888_101_fu_21735_p2 ^ Range2_all_ones_99_reg_41968);

assign deleted_zeros_99_fu_21886_p2 = (or_ln888_102_fu_21880_p2 ^ Range2_all_ones_100_reg_41997);

assign deleted_zeros_fu_18989_p2 = (or_ln888_fu_18984_p2 ^ Range2_all_ones_reg_41357);

assign lhs_100_fu_30378_p3 = ((or_ln302_109_fu_30356_p2[0:0] == 1'b1) ? select_ln302_219_fu_30362_p3 : select_ln350_109_fu_30370_p3);

assign lhs_101_fu_30480_p3 = ((or_ln302_110_fu_30458_p2[0:0] == 1'b1) ? select_ln302_221_fu_30464_p3 : select_ln350_110_fu_30472_p3);

assign lhs_102_fu_30582_p3 = ((or_ln302_111_fu_30560_p2[0:0] == 1'b1) ? select_ln302_223_fu_30566_p3 : select_ln350_111_fu_30574_p3);

assign lhs_103_fu_30684_p3 = ((or_ln302_112_fu_30662_p2[0:0] == 1'b1) ? select_ln302_225_fu_30668_p3 : select_ln350_112_fu_30676_p3);

assign lhs_104_fu_30786_p3 = ((or_ln302_113_fu_30764_p2[0:0] == 1'b1) ? select_ln302_227_fu_30770_p3 : select_ln350_113_fu_30778_p3);

assign lhs_105_fu_30888_p3 = ((or_ln302_114_fu_30866_p2[0:0] == 1'b1) ? select_ln302_229_fu_30872_p3 : select_ln350_114_fu_30880_p3);

assign lhs_106_fu_30990_p3 = ((or_ln302_115_fu_30968_p2[0:0] == 1'b1) ? select_ln302_231_fu_30974_p3 : select_ln350_115_fu_30982_p3);

assign lhs_107_fu_34768_p3 = ((or_ln302_116_fu_34748_p2[0:0] == 1'b1) ? select_ln302_233_fu_34754_p3 : select_ln350_116_fu_34761_p3);

assign lhs_108_fu_34826_p3 = ((or_ln302_117_fu_34806_p2[0:0] == 1'b1) ? select_ln302_235_fu_34812_p3 : select_ln350_117_fu_34819_p3);

assign lhs_109_fu_34884_p3 = ((or_ln302_118_fu_34864_p2[0:0] == 1'b1) ? select_ln302_237_fu_34870_p3 : select_ln350_118_fu_34877_p3);

assign lhs_110_fu_34942_p3 = ((or_ln302_119_fu_34922_p2[0:0] == 1'b1) ? select_ln302_239_fu_34928_p3 : select_ln350_119_fu_34935_p3);

assign lhs_111_fu_35000_p3 = ((or_ln302_120_fu_34980_p2[0:0] == 1'b1) ? select_ln302_241_fu_34986_p3 : select_ln350_120_fu_34993_p3);

assign lhs_112_fu_35058_p3 = ((or_ln302_121_fu_35038_p2[0:0] == 1'b1) ? select_ln302_243_fu_35044_p3 : select_ln350_121_fu_35051_p3);

assign lhs_113_fu_35116_p3 = ((or_ln302_122_fu_35096_p2[0:0] == 1'b1) ? select_ln302_245_fu_35102_p3 : select_ln350_122_fu_35109_p3);

assign lhs_114_fu_35174_p3 = ((or_ln302_123_fu_35154_p2[0:0] == 1'b1) ? select_ln302_247_fu_35160_p3 : select_ln350_123_fu_35167_p3);

assign lhs_115_fu_35232_p3 = ((or_ln302_124_fu_35212_p2[0:0] == 1'b1) ? select_ln302_249_fu_35218_p3 : select_ln350_124_fu_35225_p3);

assign lhs_116_fu_35334_p3 = ((or_ln302_125_fu_35312_p2[0:0] == 1'b1) ? select_ln302_251_fu_35318_p3 : select_ln350_125_fu_35326_p3);

assign lhs_117_fu_35436_p3 = ((or_ln302_126_fu_35414_p2[0:0] == 1'b1) ? select_ln302_253_fu_35420_p3 : select_ln350_126_fu_35428_p3);

assign lhs_118_fu_35538_p3 = ((or_ln302_127_fu_35516_p2[0:0] == 1'b1) ? select_ln302_255_fu_35522_p3 : select_ln350_127_fu_35530_p3);

assign lhs_119_fu_35640_p3 = ((or_ln302_128_fu_35618_p2[0:0] == 1'b1) ? select_ln302_257_fu_35624_p3 : select_ln350_128_fu_35632_p3);

assign lhs_120_fu_35742_p3 = ((or_ln302_129_fu_35720_p2[0:0] == 1'b1) ? select_ln302_259_fu_35726_p3 : select_ln350_129_fu_35734_p3);

assign lhs_121_fu_35844_p3 = ((or_ln302_130_fu_35822_p2[0:0] == 1'b1) ? select_ln302_261_fu_35828_p3 : select_ln350_130_fu_35836_p3);

assign lhs_122_fu_35946_p3 = ((or_ln302_131_fu_35924_p2[0:0] == 1'b1) ? select_ln302_263_fu_35930_p3 : select_ln350_131_fu_35938_p3);

assign lhs_123_fu_36048_p3 = ((or_ln302_132_fu_36026_p2[0:0] == 1'b1) ? select_ln302_265_fu_36032_p3 : select_ln350_132_fu_36040_p3);

assign lhs_124_fu_36150_p3 = ((or_ln302_133_fu_36128_p2[0:0] == 1'b1) ? select_ln302_267_fu_36134_p3 : select_ln350_133_fu_36142_p3);

assign lhs_125_fu_36252_p3 = ((or_ln302_134_fu_36230_p2[0:0] == 1'b1) ? select_ln302_269_fu_36236_p3 : select_ln350_134_fu_36244_p3);

assign lhs_126_fu_36354_p3 = ((or_ln302_135_fu_36332_p2[0:0] == 1'b1) ? select_ln302_271_fu_36338_p3 : select_ln350_135_fu_36346_p3);

assign lhs_127_fu_36456_p3 = ((or_ln302_136_fu_36434_p2[0:0] == 1'b1) ? select_ln302_273_fu_36440_p3 : select_ln350_136_fu_36448_p3);

assign lhs_128_fu_36558_p3 = ((or_ln302_137_fu_36536_p2[0:0] == 1'b1) ? select_ln302_275_fu_36542_p3 : select_ln350_137_fu_36550_p3);

assign lhs_129_fu_36660_p3 = ((or_ln302_138_fu_36638_p2[0:0] == 1'b1) ? select_ln302_277_fu_36644_p3 : select_ln350_138_fu_36652_p3);

assign lhs_130_fu_36762_p3 = ((or_ln302_139_fu_36740_p2[0:0] == 1'b1) ? select_ln302_279_fu_36746_p3 : select_ln350_139_fu_36754_p3);

assign lhs_131_fu_36864_p3 = ((or_ln302_140_fu_36842_p2[0:0] == 1'b1) ? select_ln302_281_fu_36848_p3 : select_ln350_140_fu_36856_p3);

assign lhs_132_fu_36966_p3 = ((or_ln302_141_fu_36944_p2[0:0] == 1'b1) ? select_ln302_283_fu_36950_p3 : select_ln350_141_fu_36958_p3);

assign lhs_133_fu_37068_p3 = ((or_ln302_142_fu_37046_p2[0:0] == 1'b1) ? select_ln302_285_fu_37052_p3 : select_ln350_142_fu_37060_p3);

assign lhs_134_fu_39494_p3 = ((or_ln302_143_fu_39472_p2[0:0] == 1'b1) ? select_ln302_287_fu_39478_p3 : select_ln350_143_fu_39486_p3);

assign lhs_135_fu_39594_p3 = ((or_ln302_144_fu_39572_p2[0:0] == 1'b1) ? select_ln302_289_fu_39578_p3 : select_ln350_144_fu_39586_p3);

assign lhs_136_fu_39694_p3 = ((or_ln302_145_fu_39672_p2[0:0] == 1'b1) ? select_ln302_291_fu_39678_p3 : select_ln350_145_fu_39686_p3);

assign lhs_137_fu_39794_p3 = ((or_ln302_146_fu_39772_p2[0:0] == 1'b1) ? select_ln302_293_fu_39778_p3 : select_ln350_146_fu_39786_p3);

assign lhs_138_fu_39894_p3 = ((or_ln302_147_fu_39872_p2[0:0] == 1'b1) ? select_ln302_295_fu_39878_p3 : select_ln350_147_fu_39886_p3);

assign lhs_139_fu_39994_p3 = ((or_ln302_148_fu_39972_p2[0:0] == 1'b1) ? select_ln302_297_fu_39978_p3 : select_ln350_148_fu_39986_p3);

assign lhs_140_fu_40094_p3 = ((or_ln302_149_fu_40072_p2[0:0] == 1'b1) ? select_ln302_299_fu_40078_p3 : select_ln350_149_fu_40086_p3);

assign lhs_141_fu_40194_p3 = ((or_ln302_150_fu_40172_p2[0:0] == 1'b1) ? select_ln302_301_fu_40178_p3 : select_ln350_150_fu_40186_p3);

assign lhs_142_fu_40294_p3 = ((or_ln302_151_fu_40272_p2[0:0] == 1'b1) ? select_ln302_303_fu_40278_p3 : select_ln350_151_fu_40286_p3);

assign lhs_72_fu_23810_p3 = ((or_ln302_81_fu_23788_p2[0:0] == 1'b1) ? select_ln302_163_fu_23794_p3 : select_ln350_81_fu_23802_p3);

assign lhs_73_fu_23908_p3 = ((or_ln302_82_fu_23886_p2[0:0] == 1'b1) ? select_ln302_165_fu_23892_p3 : select_ln350_82_fu_23900_p3);

assign lhs_74_fu_24006_p3 = ((or_ln302_83_fu_23984_p2[0:0] == 1'b1) ? select_ln302_167_fu_23990_p3 : select_ln350_83_fu_23998_p3);

assign lhs_75_fu_24104_p3 = ((or_ln302_84_fu_24082_p2[0:0] == 1'b1) ? select_ln302_169_fu_24088_p3 : select_ln350_84_fu_24096_p3);

assign lhs_76_fu_24202_p3 = ((or_ln302_85_fu_24180_p2[0:0] == 1'b1) ? select_ln302_171_fu_24186_p3 : select_ln350_85_fu_24194_p3);

assign lhs_77_fu_24300_p3 = ((or_ln302_86_fu_24278_p2[0:0] == 1'b1) ? select_ln302_173_fu_24284_p3 : select_ln350_86_fu_24292_p3);

assign lhs_78_fu_24398_p3 = ((or_ln302_87_fu_24376_p2[0:0] == 1'b1) ? select_ln302_175_fu_24382_p3 : select_ln350_87_fu_24390_p3);

assign lhs_79_fu_24496_p3 = ((or_ln302_88_fu_24474_p2[0:0] == 1'b1) ? select_ln302_177_fu_24480_p3 : select_ln350_88_fu_24488_p3);

assign lhs_80_fu_24598_p3 = ((or_ln302_89_fu_24576_p2[0:0] == 1'b1) ? select_ln302_179_fu_24582_p3 : select_ln350_89_fu_24590_p3);

assign lhs_81_fu_24700_p3 = ((or_ln302_90_fu_24678_p2[0:0] == 1'b1) ? select_ln302_181_fu_24684_p3 : select_ln350_90_fu_24692_p3);

assign lhs_82_fu_24802_p3 = ((or_ln302_91_fu_24780_p2[0:0] == 1'b1) ? select_ln302_183_fu_24786_p3 : select_ln350_91_fu_24794_p3);

assign lhs_83_fu_24904_p3 = ((or_ln302_92_fu_24882_p2[0:0] == 1'b1) ? select_ln302_185_fu_24888_p3 : select_ln350_92_fu_24896_p3);

assign lhs_84_fu_25006_p3 = ((or_ln302_93_fu_24984_p2[0:0] == 1'b1) ? select_ln302_187_fu_24990_p3 : select_ln350_93_fu_24998_p3);

assign lhs_85_fu_25108_p3 = ((or_ln302_94_fu_25086_p2[0:0] == 1'b1) ? select_ln302_189_fu_25092_p3 : select_ln350_94_fu_25100_p3);

assign lhs_86_fu_25210_p3 = ((or_ln302_95_fu_25188_p2[0:0] == 1'b1) ? select_ln302_191_fu_25194_p3 : select_ln350_95_fu_25202_p3);

assign lhs_87_fu_25312_p3 = ((or_ln302_96_fu_25290_p2[0:0] == 1'b1) ? select_ln302_193_fu_25296_p3 : select_ln350_96_fu_25304_p3);

assign lhs_88_fu_25414_p3 = ((or_ln302_97_fu_25392_p2[0:0] == 1'b1) ? select_ln302_195_fu_25398_p3 : select_ln350_97_fu_25406_p3);

assign lhs_89_fu_29274_p3 = ((or_ln302_98_fu_29252_p2[0:0] == 1'b1) ? select_ln302_197_fu_29258_p3 : select_ln350_98_fu_29266_p3);

assign lhs_90_fu_29374_p3 = ((or_ln302_99_fu_29352_p2[0:0] == 1'b1) ? select_ln302_199_fu_29358_p3 : select_ln350_99_fu_29366_p3);

assign lhs_91_fu_29474_p3 = ((or_ln302_100_fu_29452_p2[0:0] == 1'b1) ? select_ln302_201_fu_29458_p3 : select_ln350_100_fu_29466_p3);

assign lhs_92_fu_29572_p3 = ((or_ln302_101_fu_29550_p2[0:0] == 1'b1) ? select_ln302_203_fu_29556_p3 : select_ln350_101_fu_29564_p3);

assign lhs_93_fu_29672_p3 = ((or_ln302_102_fu_29650_p2[0:0] == 1'b1) ? select_ln302_205_fu_29656_p3 : select_ln350_102_fu_29664_p3);

assign lhs_94_fu_29772_p3 = ((or_ln302_103_fu_29750_p2[0:0] == 1'b1) ? select_ln302_207_fu_29756_p3 : select_ln350_103_fu_29764_p3);

assign lhs_95_fu_29872_p3 = ((or_ln302_104_fu_29850_p2[0:0] == 1'b1) ? select_ln302_209_fu_29856_p3 : select_ln350_104_fu_29864_p3);

assign lhs_96_fu_29972_p3 = ((or_ln302_105_fu_29950_p2[0:0] == 1'b1) ? select_ln302_211_fu_29956_p3 : select_ln350_105_fu_29964_p3);

assign lhs_97_fu_30072_p3 = ((or_ln302_106_fu_30050_p2[0:0] == 1'b1) ? select_ln302_213_fu_30056_p3 : select_ln350_106_fu_30064_p3);

assign lhs_98_fu_30174_p3 = ((or_ln302_107_fu_30152_p2[0:0] == 1'b1) ? select_ln302_215_fu_30158_p3 : select_ln350_107_fu_30166_p3);

assign lhs_99_fu_30276_p3 = ((or_ln302_108_fu_30254_p2[0:0] == 1'b1) ? select_ln302_217_fu_30260_p3 : select_ln350_108_fu_30268_p3);

assign lhs_fu_23712_p3 = ((or_ln302_fu_23690_p2[0:0] == 1'b1) ? select_ln302_fu_23696_p3 : select_ln350_fu_23704_p3);

assign or_ln302_100_fu_29452_p2 = (xor_ln302_202_fu_29446_p2 | overflow_262_fu_29422_p2);

assign or_ln302_101_fu_29550_p2 = (xor_ln302_204_fu_29544_p2 | overflow_263_fu_29520_p2);

assign or_ln302_102_fu_29650_p2 = (xor_ln302_206_fu_29644_p2 | overflow_264_fu_29620_p2);

assign or_ln302_103_fu_29750_p2 = (xor_ln302_208_fu_29744_p2 | overflow_265_fu_29720_p2);

assign or_ln302_104_fu_29850_p2 = (xor_ln302_210_fu_29844_p2 | overflow_266_fu_29820_p2);

assign or_ln302_105_fu_29950_p2 = (xor_ln302_212_fu_29944_p2 | overflow_267_fu_29920_p2);

assign or_ln302_106_fu_30050_p2 = (xor_ln302_214_fu_30044_p2 | overflow_268_fu_30020_p2);

assign or_ln302_107_fu_30152_p2 = (xor_ln302_216_fu_30146_p2 | overflow_269_fu_30122_p2);

assign or_ln302_108_fu_30254_p2 = (xor_ln302_218_fu_30248_p2 | overflow_270_fu_30224_p2);

assign or_ln302_109_fu_30356_p2 = (xor_ln302_220_fu_30350_p2 | overflow_271_fu_30326_p2);

assign or_ln302_110_fu_30458_p2 = (xor_ln302_222_fu_30452_p2 | overflow_272_fu_30428_p2);

assign or_ln302_111_fu_30560_p2 = (xor_ln302_224_fu_30554_p2 | overflow_273_fu_30530_p2);

assign or_ln302_112_fu_30662_p2 = (xor_ln302_226_fu_30656_p2 | overflow_274_fu_30632_p2);

assign or_ln302_113_fu_30764_p2 = (xor_ln302_228_fu_30758_p2 | overflow_275_fu_30734_p2);

assign or_ln302_114_fu_30866_p2 = (xor_ln302_230_fu_30860_p2 | overflow_276_fu_30836_p2);

assign or_ln302_115_fu_30968_p2 = (xor_ln302_232_fu_30962_p2 | overflow_277_fu_30938_p2);

assign or_ln302_116_fu_34748_p2 = (xor_ln302_234_fu_34742_p2 | overflow_278_fu_34723_p2);

assign or_ln302_117_fu_34806_p2 = (xor_ln302_236_fu_34800_p2 | overflow_279_fu_34781_p2);

assign or_ln302_118_fu_34864_p2 = (xor_ln302_238_fu_34858_p2 | overflow_280_fu_34839_p2);

assign or_ln302_119_fu_34922_p2 = (xor_ln302_240_fu_34916_p2 | overflow_281_fu_34897_p2);

assign or_ln302_120_fu_34980_p2 = (xor_ln302_242_fu_34974_p2 | overflow_282_fu_34955_p2);

assign or_ln302_121_fu_35038_p2 = (xor_ln302_244_fu_35032_p2 | overflow_283_fu_35013_p2);

assign or_ln302_122_fu_35096_p2 = (xor_ln302_246_fu_35090_p2 | overflow_284_fu_35071_p2);

assign or_ln302_123_fu_35154_p2 = (xor_ln302_248_fu_35148_p2 | overflow_285_fu_35129_p2);

assign or_ln302_124_fu_35212_p2 = (xor_ln302_250_fu_35206_p2 | overflow_286_fu_35187_p2);

assign or_ln302_125_fu_35312_p2 = (xor_ln302_252_fu_35306_p2 | overflow_287_fu_35282_p2);

assign or_ln302_126_fu_35414_p2 = (xor_ln302_254_fu_35408_p2 | overflow_288_fu_35384_p2);

assign or_ln302_127_fu_35516_p2 = (xor_ln302_256_fu_35510_p2 | overflow_289_fu_35486_p2);

assign or_ln302_128_fu_35618_p2 = (xor_ln302_258_fu_35612_p2 | overflow_290_fu_35588_p2);

assign or_ln302_129_fu_35720_p2 = (xor_ln302_260_fu_35714_p2 | overflow_291_fu_35690_p2);

assign or_ln302_130_fu_35822_p2 = (xor_ln302_262_fu_35816_p2 | overflow_292_fu_35792_p2);

assign or_ln302_131_fu_35924_p2 = (xor_ln302_264_fu_35918_p2 | overflow_293_fu_35894_p2);

assign or_ln302_132_fu_36026_p2 = (xor_ln302_266_fu_36020_p2 | overflow_294_fu_35996_p2);

assign or_ln302_133_fu_36128_p2 = (xor_ln302_268_fu_36122_p2 | overflow_295_fu_36098_p2);

assign or_ln302_134_fu_36230_p2 = (xor_ln302_270_fu_36224_p2 | overflow_296_fu_36200_p2);

assign or_ln302_135_fu_36332_p2 = (xor_ln302_272_fu_36326_p2 | overflow_297_fu_36302_p2);

assign or_ln302_136_fu_36434_p2 = (xor_ln302_274_fu_36428_p2 | overflow_298_fu_36404_p2);

assign or_ln302_137_fu_36536_p2 = (xor_ln302_276_fu_36530_p2 | overflow_299_fu_36506_p2);

assign or_ln302_138_fu_36638_p2 = (xor_ln302_278_fu_36632_p2 | overflow_300_fu_36608_p2);

assign or_ln302_139_fu_36740_p2 = (xor_ln302_280_fu_36734_p2 | overflow_301_fu_36710_p2);

assign or_ln302_140_fu_36842_p2 = (xor_ln302_282_fu_36836_p2 | overflow_302_fu_36812_p2);

assign or_ln302_141_fu_36944_p2 = (xor_ln302_284_fu_36938_p2 | overflow_303_fu_36914_p2);

assign or_ln302_142_fu_37046_p2 = (xor_ln302_286_fu_37040_p2 | overflow_304_fu_37016_p2);

assign or_ln302_143_fu_39472_p2 = (xor_ln302_288_fu_39466_p2 | overflow_305_fu_39442_p2);

assign or_ln302_144_fu_39572_p2 = (xor_ln302_290_fu_39566_p2 | overflow_306_fu_39542_p2);

assign or_ln302_145_fu_39672_p2 = (xor_ln302_292_fu_39666_p2 | overflow_307_fu_39642_p2);

assign or_ln302_146_fu_39772_p2 = (xor_ln302_294_fu_39766_p2 | overflow_308_fu_39742_p2);

assign or_ln302_147_fu_39872_p2 = (xor_ln302_296_fu_39866_p2 | overflow_309_fu_39842_p2);

assign or_ln302_148_fu_39972_p2 = (xor_ln302_298_fu_39966_p2 | overflow_310_fu_39942_p2);

assign or_ln302_149_fu_40072_p2 = (xor_ln302_300_fu_40066_p2 | overflow_311_fu_40042_p2);

assign or_ln302_150_fu_40172_p2 = (xor_ln302_302_fu_40166_p2 | overflow_312_fu_40142_p2);

assign or_ln302_151_fu_40272_p2 = (xor_ln302_304_fu_40266_p2 | overflow_313_fu_40242_p2);

assign or_ln302_152_fu_40374_p2 = (xor_ln302_306_fu_40368_p2 | overflow_314_fu_40344_p2);

assign or_ln302_153_fu_40476_p2 = (xor_ln302_308_fu_40470_p2 | overflow_315_fu_40446_p2);

assign or_ln302_154_fu_40578_p2 = (xor_ln302_310_fu_40572_p2 | overflow_316_fu_40548_p2);

assign or_ln302_155_fu_40680_p2 = (xor_ln302_312_fu_40674_p2 | overflow_317_fu_40650_p2);

assign or_ln302_156_fu_40782_p2 = (xor_ln302_314_fu_40776_p2 | overflow_318_fu_40752_p2);

assign or_ln302_157_fu_40884_p2 = (xor_ln302_316_fu_40878_p2 | overflow_319_fu_40854_p2);

assign or_ln302_158_fu_40986_p2 = (xor_ln302_318_fu_40980_p2 | overflow_320_fu_40956_p2);

assign or_ln302_159_fu_41088_p2 = (xor_ln302_320_fu_41082_p2 | overflow_321_fu_41058_p2);

assign or_ln302_160_fu_41190_p2 = (xor_ln302_322_fu_41184_p2 | overflow_322_fu_41160_p2);

assign or_ln302_81_fu_23788_p2 = (xor_ln302_164_fu_23782_p2 | overflow_243_fu_23758_p2);

assign or_ln302_82_fu_23886_p2 = (xor_ln302_166_fu_23880_p2 | overflow_244_fu_23856_p2);

assign or_ln302_83_fu_23984_p2 = (xor_ln302_168_fu_23978_p2 | overflow_245_fu_23954_p2);

assign or_ln302_84_fu_24082_p2 = (xor_ln302_170_fu_24076_p2 | overflow_246_fu_24052_p2);

assign or_ln302_85_fu_24180_p2 = (xor_ln302_172_fu_24174_p2 | overflow_247_fu_24150_p2);

assign or_ln302_86_fu_24278_p2 = (xor_ln302_174_fu_24272_p2 | overflow_248_fu_24248_p2);

assign or_ln302_87_fu_24376_p2 = (xor_ln302_176_fu_24370_p2 | overflow_249_fu_24346_p2);

assign or_ln302_88_fu_24474_p2 = (xor_ln302_178_fu_24468_p2 | overflow_250_fu_24444_p2);

assign or_ln302_89_fu_24576_p2 = (xor_ln302_180_fu_24570_p2 | overflow_251_fu_24546_p2);

assign or_ln302_90_fu_24678_p2 = (xor_ln302_182_fu_24672_p2 | overflow_252_fu_24648_p2);

assign or_ln302_91_fu_24780_p2 = (xor_ln302_184_fu_24774_p2 | overflow_253_fu_24750_p2);

assign or_ln302_92_fu_24882_p2 = (xor_ln302_186_fu_24876_p2 | overflow_254_fu_24852_p2);

assign or_ln302_93_fu_24984_p2 = (xor_ln302_188_fu_24978_p2 | overflow_255_fu_24954_p2);

assign or_ln302_94_fu_25086_p2 = (xor_ln302_190_fu_25080_p2 | overflow_256_fu_25056_p2);

assign or_ln302_95_fu_25188_p2 = (xor_ln302_192_fu_25182_p2 | overflow_257_fu_25158_p2);

assign or_ln302_96_fu_25290_p2 = (xor_ln302_194_fu_25284_p2 | overflow_258_fu_25260_p2);

assign or_ln302_97_fu_25392_p2 = (xor_ln302_196_fu_25386_p2 | overflow_259_fu_25362_p2);

assign or_ln302_98_fu_29252_p2 = (xor_ln302_198_fu_29246_p2 | overflow_260_fu_29222_p2);

assign or_ln302_99_fu_29352_p2 = (xor_ln302_200_fu_29346_p2 | overflow_261_fu_29322_p2);

assign or_ln302_fu_23690_p2 = (xor_ln302_162_fu_23684_p2 | overflow_242_fu_23660_p2);

assign or_ln346_100_fu_21697_p2 = (underflow_181_fu_21692_p2 | overflow_181_fu_21668_p2);

assign or_ln346_101_fu_21830_p2 = (underflow_182_fu_21817_p2 | overflow_182_fu_21793_p2);

assign or_ln346_102_fu_21967_p2 = (underflow_183_fu_21962_p2 | overflow_183_fu_21938_p2);

assign or_ln346_103_fu_22096_p2 = (underflow_184_fu_22091_p2 | overflow_184_fu_22067_p2);

assign or_ln346_104_fu_22225_p2 = (underflow_185_fu_22220_p2 | overflow_185_fu_22196_p2);

assign or_ln346_105_fu_22354_p2 = (underflow_186_fu_22349_p2 | overflow_186_fu_22325_p2);

assign or_ln346_106_fu_22483_p2 = (underflow_187_fu_22478_p2 | overflow_187_fu_22454_p2);

assign or_ln346_107_fu_25652_p2 = (underflow_188_fu_25639_p2 | overflow_188_fu_25615_p2);

assign or_ln346_108_fu_25777_p2 = (underflow_189_fu_25764_p2 | overflow_189_fu_25740_p2);

assign or_ln346_109_fu_25902_p2 = (underflow_190_fu_25889_p2 | overflow_190_fu_25865_p2);

assign or_ln346_110_fu_26027_p2 = (underflow_191_fu_26014_p2 | overflow_191_fu_25990_p2);

assign or_ln346_111_fu_26152_p2 = (underflow_192_fu_26139_p2 | overflow_192_fu_26115_p2);

assign or_ln346_112_fu_26277_p2 = (underflow_193_fu_26264_p2 | overflow_193_fu_26240_p2);

assign or_ln346_113_fu_23083_p2 = (underflow_194_fu_23077_p2 | overflow_194_fu_23053_p2);

assign or_ln346_114_fu_26419_p2 = (underflow_195_fu_26406_p2 | overflow_195_fu_26382_p2);

assign or_ln346_115_fu_26544_p2 = (underflow_196_fu_26531_p2 | overflow_196_fu_26507_p2);

assign or_ln346_116_fu_26689_p2 = (underflow_197_fu_26676_p2 | overflow_197_fu_26652_p2);

assign or_ln346_117_fu_26838_p2 = (underflow_198_fu_26825_p2 | overflow_198_fu_26801_p2);

assign or_ln346_118_fu_26987_p2 = (underflow_199_fu_26974_p2 | overflow_199_fu_26950_p2);

assign or_ln346_119_fu_27136_p2 = (underflow_200_fu_27123_p2 | overflow_200_fu_27099_p2);

assign or_ln346_120_fu_27285_p2 = (underflow_201_fu_27272_p2 | overflow_201_fu_27248_p2);

assign or_ln346_121_fu_27434_p2 = (underflow_202_fu_27421_p2 | overflow_202_fu_27397_p2);

assign or_ln346_122_fu_27583_p2 = (underflow_203_fu_27570_p2 | overflow_203_fu_27546_p2);

assign or_ln346_123_fu_27732_p2 = (underflow_204_fu_27719_p2 | overflow_204_fu_27695_p2);

assign or_ln346_124_fu_27881_p2 = (underflow_205_fu_27868_p2 | overflow_205_fu_27844_p2);

assign or_ln346_125_fu_28111_p2 = (underflow_206_fu_28105_p2 | overflow_206_fu_28081_p2);

assign or_ln346_126_fu_31450_p2 = (underflow_207_fu_31437_p2 | overflow_207_fu_31413_p2);

assign or_ln346_127_fu_31575_p2 = (underflow_208_fu_31562_p2 | overflow_208_fu_31538_p2);

assign or_ln346_128_fu_31700_p2 = (underflow_209_fu_31687_p2 | overflow_209_fu_31663_p2);

assign or_ln346_129_fu_31825_p2 = (underflow_210_fu_31812_p2 | overflow_210_fu_31788_p2);

assign or_ln346_130_fu_31950_p2 = (underflow_211_fu_31937_p2 | overflow_211_fu_31913_p2);

assign or_ln346_131_fu_32075_p2 = (underflow_212_fu_32062_p2 | overflow_212_fu_32038_p2);

assign or_ln346_132_fu_32200_p2 = (underflow_213_fu_32187_p2 | overflow_213_fu_32163_p2);

assign or_ln346_133_fu_32325_p2 = (underflow_214_fu_32312_p2 | overflow_214_fu_32288_p2);

assign or_ln346_134_fu_32474_p2 = (underflow_215_fu_32461_p2 | overflow_215_fu_32437_p2);

assign or_ln346_135_fu_32623_p2 = (underflow_216_fu_32610_p2 | overflow_216_fu_32586_p2);

assign or_ln346_136_fu_32772_p2 = (underflow_217_fu_32759_p2 | overflow_217_fu_32735_p2);

assign or_ln346_137_fu_32921_p2 = (underflow_218_fu_32908_p2 | overflow_218_fu_32884_p2);

assign or_ln346_138_fu_33070_p2 = (underflow_219_fu_33057_p2 | overflow_219_fu_33033_p2);

assign or_ln346_139_fu_33219_p2 = (underflow_220_fu_33206_p2 | overflow_220_fu_33182_p2);

assign or_ln346_140_fu_33368_p2 = (underflow_221_fu_33355_p2 | overflow_221_fu_33331_p2);

assign or_ln346_141_fu_33517_p2 = (underflow_222_fu_33504_p2 | overflow_222_fu_33480_p2);

assign or_ln346_142_fu_29178_p2 = (underflow_223_fu_29172_p2 | overflow_223_fu_29148_p2);

assign or_ln346_143_fu_37184_p2 = (underflow_224_fu_37171_p2 | overflow_224_fu_37147_p2);

assign or_ln346_144_fu_37308_p2 = (underflow_225_fu_37295_p2 | overflow_225_fu_37271_p2);

assign or_ln346_145_fu_37433_p2 = (underflow_226_fu_37420_p2 | overflow_226_fu_37396_p2);

assign or_ln346_146_fu_37558_p2 = (underflow_227_fu_37545_p2 | overflow_227_fu_37521_p2);

assign or_ln346_147_fu_37683_p2 = (underflow_228_fu_37670_p2 | overflow_228_fu_37646_p2);

assign or_ln346_148_fu_37808_p2 = (underflow_229_fu_37795_p2 | overflow_229_fu_37771_p2);

assign or_ln346_149_fu_37933_p2 = (underflow_230_fu_37920_p2 | overflow_230_fu_37896_p2);

assign or_ln346_150_fu_38058_p2 = (underflow_231_fu_38045_p2 | overflow_231_fu_38021_p2);

assign or_ln346_151_fu_38183_p2 = (underflow_232_fu_38170_p2 | overflow_232_fu_38146_p2);

assign or_ln346_152_fu_38328_p2 = (underflow_233_fu_38315_p2 | overflow_233_fu_38291_p2);

assign or_ln346_153_fu_38477_p2 = (underflow_234_fu_38464_p2 | overflow_234_fu_38440_p2);

assign or_ln346_154_fu_38626_p2 = (underflow_235_fu_38613_p2 | overflow_235_fu_38589_p2);

assign or_ln346_155_fu_38775_p2 = (underflow_236_fu_38762_p2 | overflow_236_fu_38738_p2);

assign or_ln346_156_fu_38924_p2 = (underflow_237_fu_38911_p2 | overflow_237_fu_38887_p2);

assign or_ln346_157_fu_39073_p2 = (underflow_238_fu_39060_p2 | overflow_238_fu_39036_p2);

assign or_ln346_158_fu_39222_p2 = (underflow_239_fu_39209_p2 | overflow_239_fu_39185_p2);

assign or_ln346_159_fu_34670_p2 = (underflow_240_fu_34664_p2 | overflow_240_fu_34640_p2);

assign or_ln346_160_fu_39388_p2 = (underflow_241_fu_39375_p2 | overflow_241_fu_39351_p2);

assign or_ln346_81_fu_19202_p2 = (underflow_162_fu_19189_p2 | overflow_162_fu_19165_p2);

assign or_ln346_82_fu_19327_p2 = (underflow_163_fu_19314_p2 | overflow_163_fu_19290_p2);

assign or_ln346_83_fu_19452_p2 = (underflow_164_fu_19439_p2 | overflow_164_fu_19415_p2);

assign or_ln346_84_fu_19577_p2 = (underflow_165_fu_19564_p2 | overflow_165_fu_19540_p2);

assign or_ln346_85_fu_19702_p2 = (underflow_166_fu_19689_p2 | overflow_166_fu_19665_p2);

assign or_ln346_86_fu_19827_p2 = (underflow_167_fu_19814_p2 | overflow_167_fu_19790_p2);

assign or_ln346_87_fu_19952_p2 = (underflow_168_fu_19939_p2 | overflow_168_fu_19915_p2);

assign or_ln346_88_fu_20077_p2 = (underflow_169_fu_20064_p2 | overflow_169_fu_20040_p2);

assign or_ln346_89_fu_20226_p2 = (underflow_170_fu_20213_p2 | overflow_170_fu_20189_p2);

assign or_ln346_90_fu_20375_p2 = (underflow_171_fu_20362_p2 | overflow_171_fu_20338_p2);

assign or_ln346_91_fu_20524_p2 = (underflow_172_fu_20511_p2 | overflow_172_fu_20487_p2);

assign or_ln346_92_fu_20673_p2 = (underflow_173_fu_20660_p2 | overflow_173_fu_20636_p2);

assign or_ln346_93_fu_20822_p2 = (underflow_174_fu_20809_p2 | overflow_174_fu_20785_p2);

assign or_ln346_94_fu_18301_p2 = (underflow_175_fu_18295_p2 | overflow_175_fu_18271_p2);

assign or_ln346_95_fu_20988_p2 = (underflow_176_fu_20975_p2 | overflow_176_fu_20951_p2);

assign or_ln346_96_fu_21137_p2 = (underflow_177_fu_21124_p2 | overflow_177_fu_21100_p2);

assign or_ln346_97_fu_21286_p2 = (underflow_178_fu_21273_p2 | overflow_178_fu_21249_p2);

assign or_ln346_98_fu_21431_p2 = (underflow_179_fu_21418_p2 | overflow_179_fu_21394_p2);

assign or_ln346_99_fu_21568_p2 = (underflow_180_fu_21563_p2 | overflow_180_fu_21539_p2);

assign or_ln346_fu_19077_p2 = (underflow_fu_19064_p2 | overflow_fu_19040_p2);

assign or_ln888_100_fu_21610_p2 = (xor_ln888_198_fu_21605_p2 | p_Result_464_fu_21586_p3);

assign or_ln888_101_fu_21735_p2 = (xor_ln888_200_fu_21730_p2 | p_Result_467_fu_21711_p3);

assign or_ln888_102_fu_21880_p2 = (xor_ln888_202_fu_21875_p2 | p_Result_470_fu_21856_p3);

assign or_ln888_103_fu_22009_p2 = (xor_ln888_204_fu_22004_p2 | p_Result_473_fu_21985_p3);

assign or_ln888_104_fu_22138_p2 = (xor_ln888_206_fu_22133_p2 | p_Result_476_fu_22114_p3);

assign or_ln888_105_fu_22267_p2 = (xor_ln888_208_fu_22262_p2 | p_Result_479_fu_22243_p3);

assign or_ln888_106_fu_22396_p2 = (xor_ln888_210_fu_22391_p2 | p_Result_482_fu_22372_p3);

assign or_ln888_107_fu_25559_p2 = (xor_ln888_212_fu_25554_p2 | p_Result_485_reg_42269);

assign or_ln888_108_fu_25684_p2 = (xor_ln888_214_fu_25679_p2 | p_Result_488_reg_42300);

assign or_ln888_109_fu_25809_p2 = (xor_ln888_216_fu_25804_p2 | p_Result_491_reg_42331);

assign or_ln888_110_fu_25934_p2 = (xor_ln888_218_fu_25929_p2 | p_Result_494_reg_42362);

assign or_ln888_111_fu_26059_p2 = (xor_ln888_220_fu_26054_p2 | p_Result_497_reg_42393);

assign or_ln888_112_fu_26184_p2 = (xor_ln888_222_fu_26179_p2 | p_Result_500_reg_42424);

assign or_ln888_113_fu_22991_p2 = (xor_ln888_224_fu_22985_p2 | p_Result_503_fu_22957_p3);

assign or_ln888_114_fu_26326_p2 = (xor_ln888_226_fu_26321_p2 | p_Result_506_reg_42470);

assign or_ln888_115_fu_26451_p2 = (xor_ln888_228_fu_26446_p2 | p_Result_509_reg_42501);

assign or_ln888_116_fu_26594_p2 = (xor_ln888_230_fu_26589_p2 | p_Result_512_fu_26570_p3);

assign or_ln888_117_fu_26743_p2 = (xor_ln888_232_fu_26738_p2 | p_Result_515_fu_26719_p3);

assign or_ln888_118_fu_26892_p2 = (xor_ln888_234_fu_26887_p2 | p_Result_518_fu_26868_p3);

assign or_ln888_119_fu_27041_p2 = (xor_ln888_236_fu_27036_p2 | p_Result_521_fu_27017_p3);

assign or_ln888_120_fu_27190_p2 = (xor_ln888_238_fu_27185_p2 | p_Result_524_fu_27166_p3);

assign or_ln888_121_fu_27339_p2 = (xor_ln888_240_fu_27334_p2 | p_Result_527_fu_27315_p3);

assign or_ln888_122_fu_27488_p2 = (xor_ln888_242_fu_27483_p2 | p_Result_530_fu_27464_p3);

assign or_ln888_123_fu_27637_p2 = (xor_ln888_244_fu_27632_p2 | p_Result_533_fu_27613_p3);

assign or_ln888_124_fu_27786_p2 = (xor_ln888_246_fu_27781_p2 | p_Result_536_fu_27762_p3);

assign or_ln888_125_fu_28019_p2 = (xor_ln888_248_fu_28013_p2 | p_Result_539_fu_27985_p3);

assign or_ln888_126_fu_31357_p2 = (xor_ln888_250_fu_31352_p2 | p_Result_542_reg_42862);

assign or_ln888_127_fu_31482_p2 = (xor_ln888_252_fu_31477_p2 | p_Result_545_reg_42893);

assign or_ln888_128_fu_31607_p2 = (xor_ln888_254_fu_31602_p2 | p_Result_548_reg_42924);

assign or_ln888_129_fu_31732_p2 = (xor_ln888_256_fu_31727_p2 | p_Result_551_reg_42955);

assign or_ln888_130_fu_31857_p2 = (xor_ln888_258_fu_31852_p2 | p_Result_554_reg_42986);

assign or_ln888_131_fu_31982_p2 = (xor_ln888_260_fu_31977_p2 | p_Result_557_reg_43017);

assign or_ln888_132_fu_32107_p2 = (xor_ln888_262_fu_32102_p2 | p_Result_560_reg_43048);

assign or_ln888_133_fu_32232_p2 = (xor_ln888_264_fu_32227_p2 | p_Result_563_reg_43079);

assign or_ln888_134_fu_32379_p2 = (xor_ln888_266_fu_32374_p2 | p_Result_566_fu_32355_p3);

assign or_ln888_135_fu_32528_p2 = (xor_ln888_268_fu_32523_p2 | p_Result_569_fu_32504_p3);

assign or_ln888_136_fu_32677_p2 = (xor_ln888_270_fu_32672_p2 | p_Result_572_fu_32653_p3);

assign or_ln888_137_fu_32826_p2 = (xor_ln888_272_fu_32821_p2 | p_Result_575_fu_32802_p3);

assign or_ln888_138_fu_32975_p2 = (xor_ln888_274_fu_32970_p2 | p_Result_578_fu_32951_p3);

assign or_ln888_139_fu_33124_p2 = (xor_ln888_276_fu_33119_p2 | p_Result_581_fu_33100_p3);

assign or_ln888_140_fu_33273_p2 = (xor_ln888_278_fu_33268_p2 | p_Result_584_fu_33249_p3);

assign or_ln888_141_fu_33422_p2 = (xor_ln888_280_fu_33417_p2 | p_Result_587_fu_33398_p3);

assign or_ln888_142_fu_29086_p2 = (xor_ln888_282_fu_29080_p2 | p_Result_590_fu_29052_p3);

assign or_ln888_143_fu_37091_p2 = (xor_ln888_284_fu_37086_p2 | p_Result_593_reg_43537);

assign or_ln888_144_fu_37215_p2 = (xor_ln888_286_fu_37210_p2 | p_Result_596_reg_43568);

assign or_ln888_145_fu_37340_p2 = (xor_ln888_288_fu_37335_p2 | p_Result_599_reg_43599);

assign or_ln888_146_fu_37465_p2 = (xor_ln888_290_fu_37460_p2 | p_Result_602_reg_43630);

assign or_ln888_147_fu_37590_p2 = (xor_ln888_292_fu_37585_p2 | p_Result_605_reg_43661);

assign or_ln888_148_fu_37715_p2 = (xor_ln888_294_fu_37710_p2 | p_Result_608_reg_43692);

assign or_ln888_149_fu_37840_p2 = (xor_ln888_296_fu_37835_p2 | p_Result_611_reg_43723);

assign or_ln888_150_fu_37965_p2 = (xor_ln888_298_fu_37960_p2 | p_Result_614_reg_43754);

assign or_ln888_151_fu_38090_p2 = (xor_ln888_300_fu_38085_p2 | p_Result_617_reg_43785);

assign or_ln888_152_fu_38233_p2 = (xor_ln888_302_fu_38228_p2 | p_Result_620_fu_38209_p3);

assign or_ln888_153_fu_38382_p2 = (xor_ln888_304_fu_38377_p2 | p_Result_623_fu_38358_p3);

assign or_ln888_154_fu_38531_p2 = (xor_ln888_306_fu_38526_p2 | p_Result_626_fu_38507_p3);

assign or_ln888_155_fu_38680_p2 = (xor_ln888_308_fu_38675_p2 | p_Result_629_fu_38656_p3);

assign or_ln888_156_fu_38829_p2 = (xor_ln888_310_fu_38824_p2 | p_Result_632_fu_38805_p3);

assign or_ln888_157_fu_38978_p2 = (xor_ln888_312_fu_38973_p2 | p_Result_635_fu_38954_p3);

assign or_ln888_158_fu_39127_p2 = (xor_ln888_314_fu_39122_p2 | p_Result_638_fu_39103_p3);

assign or_ln888_159_fu_34578_p2 = (xor_ln888_316_fu_34572_p2 | p_Result_641_fu_34544_p3);

assign or_ln888_160_fu_39293_p2 = (xor_ln888_318_fu_39288_p2 | p_Result_644_fu_39269_p3);

assign or_ln888_81_fu_19109_p2 = (xor_ln888_160_fu_19104_p2 | p_Result_407_reg_41381);

assign or_ln888_82_fu_19234_p2 = (xor_ln888_162_fu_19229_p2 | p_Result_410_reg_41412);

assign or_ln888_83_fu_19359_p2 = (xor_ln888_164_fu_19354_p2 | p_Result_413_reg_41443);

assign or_ln888_84_fu_19484_p2 = (xor_ln888_166_fu_19479_p2 | p_Result_416_reg_41474);

assign or_ln888_85_fu_19609_p2 = (xor_ln888_168_fu_19604_p2 | p_Result_419_reg_41505);

assign or_ln888_86_fu_19734_p2 = (xor_ln888_170_fu_19729_p2 | p_Result_422_reg_41536);

assign or_ln888_87_fu_19859_p2 = (xor_ln888_172_fu_19854_p2 | p_Result_425_reg_41567);

assign or_ln888_88_fu_19984_p2 = (xor_ln888_174_fu_19979_p2 | p_Result_428_reg_41598);

assign or_ln888_89_fu_20131_p2 = (xor_ln888_176_fu_20126_p2 | p_Result_431_fu_20107_p3);

assign or_ln888_90_fu_20280_p2 = (xor_ln888_178_fu_20275_p2 | p_Result_434_fu_20256_p3);

assign or_ln888_91_fu_20429_p2 = (xor_ln888_180_fu_20424_p2 | p_Result_437_fu_20405_p3);

assign or_ln888_92_fu_20578_p2 = (xor_ln888_182_fu_20573_p2 | p_Result_440_fu_20554_p3);

assign or_ln888_93_fu_20727_p2 = (xor_ln888_184_fu_20722_p2 | p_Result_443_fu_20703_p3);

assign or_ln888_94_fu_18209_p2 = (xor_ln888_186_fu_18203_p2 | p_Result_446_fu_18175_p3);

assign or_ln888_95_fu_20893_p2 = (xor_ln888_188_fu_20888_p2 | p_Result_449_fu_20869_p3);

assign or_ln888_96_fu_21042_p2 = (xor_ln888_190_fu_21037_p2 | p_Result_452_fu_21018_p3);

assign or_ln888_97_fu_21191_p2 = (xor_ln888_192_fu_21186_p2 | p_Result_455_fu_21167_p3);

assign or_ln888_98_fu_21336_p2 = (xor_ln888_194_fu_21331_p2 | p_Result_458_fu_21312_p3);

assign or_ln888_99_fu_21481_p2 = (xor_ln888_196_fu_21476_p2 | p_Result_461_fu_21457_p3);

assign or_ln888_fu_18984_p2 = (xor_ln888_fu_18979_p2 | p_Result_404_reg_41350);

assign or_ln890_100_fu_21635_p2 = (xor_ln890_98_fu_21629_p2 | or_ln888_100_fu_21610_p2);

assign or_ln890_101_fu_21760_p2 = (xor_ln890_99_fu_21754_p2 | or_ln888_101_fu_21735_p2);

assign or_ln890_102_fu_21905_p2 = (xor_ln890_100_fu_21899_p2 | or_ln888_102_fu_21880_p2);

assign or_ln890_103_fu_22034_p2 = (xor_ln890_101_fu_22028_p2 | or_ln888_103_fu_22009_p2);

assign or_ln890_104_fu_22163_p2 = (xor_ln890_102_fu_22157_p2 | or_ln888_104_fu_22138_p2);

assign or_ln890_105_fu_22292_p2 = (xor_ln890_103_fu_22286_p2 | or_ln888_105_fu_22267_p2);

assign or_ln890_106_fu_22421_p2 = (xor_ln890_104_fu_22415_p2 | or_ln888_106_fu_22396_p2);

assign or_ln890_107_fu_25583_p2 = (xor_ln890_105_fu_25577_p2 | or_ln888_107_fu_25559_p2);

assign or_ln890_108_fu_25708_p2 = (xor_ln890_106_fu_25702_p2 | or_ln888_108_fu_25684_p2);

assign or_ln890_109_fu_25833_p2 = (xor_ln890_107_fu_25827_p2 | or_ln888_109_fu_25809_p2);

assign or_ln890_110_fu_25958_p2 = (xor_ln890_108_fu_25952_p2 | or_ln888_110_fu_25934_p2);

assign or_ln890_111_fu_26083_p2 = (xor_ln890_109_fu_26077_p2 | or_ln888_111_fu_26059_p2);

assign or_ln890_112_fu_26208_p2 = (xor_ln890_110_fu_26202_p2 | or_ln888_112_fu_26184_p2);

assign or_ln890_113_fu_23017_p2 = (xor_ln890_111_fu_23011_p2 | or_ln888_113_fu_22991_p2);

assign or_ln890_114_fu_26350_p2 = (xor_ln890_112_fu_26344_p2 | or_ln888_114_fu_26326_p2);

assign or_ln890_115_fu_26475_p2 = (xor_ln890_113_fu_26469_p2 | or_ln888_115_fu_26451_p2);

assign or_ln890_116_fu_26619_p2 = (xor_ln890_114_fu_26613_p2 | or_ln888_116_fu_26594_p2);

assign or_ln890_117_fu_26768_p2 = (xor_ln890_115_fu_26762_p2 | or_ln888_117_fu_26743_p2);

assign or_ln890_118_fu_26917_p2 = (xor_ln890_116_fu_26911_p2 | or_ln888_118_fu_26892_p2);

assign or_ln890_119_fu_27066_p2 = (xor_ln890_117_fu_27060_p2 | or_ln888_119_fu_27041_p2);

assign or_ln890_120_fu_27215_p2 = (xor_ln890_118_fu_27209_p2 | or_ln888_120_fu_27190_p2);

assign or_ln890_121_fu_27364_p2 = (xor_ln890_119_fu_27358_p2 | or_ln888_121_fu_27339_p2);

assign or_ln890_122_fu_27513_p2 = (xor_ln890_120_fu_27507_p2 | or_ln888_122_fu_27488_p2);

assign or_ln890_123_fu_27662_p2 = (xor_ln890_121_fu_27656_p2 | or_ln888_123_fu_27637_p2);

assign or_ln890_124_fu_27811_p2 = (xor_ln890_122_fu_27805_p2 | or_ln888_124_fu_27786_p2);

assign or_ln890_125_fu_28045_p2 = (xor_ln890_123_fu_28039_p2 | or_ln888_125_fu_28019_p2);

assign or_ln890_126_fu_31381_p2 = (xor_ln890_124_fu_31375_p2 | or_ln888_126_fu_31357_p2);

assign or_ln890_127_fu_31506_p2 = (xor_ln890_125_fu_31500_p2 | or_ln888_127_fu_31482_p2);

assign or_ln890_128_fu_31631_p2 = (xor_ln890_126_fu_31625_p2 | or_ln888_128_fu_31607_p2);

assign or_ln890_129_fu_31756_p2 = (xor_ln890_127_fu_31750_p2 | or_ln888_129_fu_31732_p2);

assign or_ln890_130_fu_31881_p2 = (xor_ln890_128_fu_31875_p2 | or_ln888_130_fu_31857_p2);

assign or_ln890_131_fu_32006_p2 = (xor_ln890_129_fu_32000_p2 | or_ln888_131_fu_31982_p2);

assign or_ln890_132_fu_32131_p2 = (xor_ln890_130_fu_32125_p2 | or_ln888_132_fu_32107_p2);

assign or_ln890_133_fu_32256_p2 = (xor_ln890_131_fu_32250_p2 | or_ln888_133_fu_32232_p2);

assign or_ln890_134_fu_32404_p2 = (xor_ln890_132_fu_32398_p2 | or_ln888_134_fu_32379_p2);

assign or_ln890_135_fu_32553_p2 = (xor_ln890_133_fu_32547_p2 | or_ln888_135_fu_32528_p2);

assign or_ln890_136_fu_32702_p2 = (xor_ln890_134_fu_32696_p2 | or_ln888_136_fu_32677_p2);

assign or_ln890_137_fu_32851_p2 = (xor_ln890_135_fu_32845_p2 | or_ln888_137_fu_32826_p2);

assign or_ln890_138_fu_33000_p2 = (xor_ln890_136_fu_32994_p2 | or_ln888_138_fu_32975_p2);

assign or_ln890_139_fu_33149_p2 = (xor_ln890_137_fu_33143_p2 | or_ln888_139_fu_33124_p2);

assign or_ln890_140_fu_33298_p2 = (xor_ln890_138_fu_33292_p2 | or_ln888_140_fu_33273_p2);

assign or_ln890_141_fu_33447_p2 = (xor_ln890_139_fu_33441_p2 | or_ln888_141_fu_33422_p2);

assign or_ln890_142_fu_29112_p2 = (xor_ln890_140_fu_29106_p2 | or_ln888_142_fu_29086_p2);

assign or_ln890_143_fu_37115_p2 = (xor_ln890_141_fu_37109_p2 | or_ln888_143_fu_37091_p2);

assign or_ln890_144_fu_37239_p2 = (xor_ln890_142_fu_37233_p2 | or_ln888_144_fu_37215_p2);

assign or_ln890_145_fu_37364_p2 = (xor_ln890_143_fu_37358_p2 | or_ln888_145_fu_37340_p2);

assign or_ln890_146_fu_37489_p2 = (xor_ln890_144_fu_37483_p2 | or_ln888_146_fu_37465_p2);

assign or_ln890_147_fu_37614_p2 = (xor_ln890_145_fu_37608_p2 | or_ln888_147_fu_37590_p2);

assign or_ln890_148_fu_37739_p2 = (xor_ln890_146_fu_37733_p2 | or_ln888_148_fu_37715_p2);

assign or_ln890_149_fu_37864_p2 = (xor_ln890_147_fu_37858_p2 | or_ln888_149_fu_37840_p2);

assign or_ln890_150_fu_37989_p2 = (xor_ln890_148_fu_37983_p2 | or_ln888_150_fu_37965_p2);

assign or_ln890_151_fu_38114_p2 = (xor_ln890_149_fu_38108_p2 | or_ln888_151_fu_38090_p2);

assign or_ln890_152_fu_38258_p2 = (xor_ln890_150_fu_38252_p2 | or_ln888_152_fu_38233_p2);

assign or_ln890_153_fu_38407_p2 = (xor_ln890_151_fu_38401_p2 | or_ln888_153_fu_38382_p2);

assign or_ln890_154_fu_38556_p2 = (xor_ln890_152_fu_38550_p2 | or_ln888_154_fu_38531_p2);

assign or_ln890_155_fu_38705_p2 = (xor_ln890_153_fu_38699_p2 | or_ln888_155_fu_38680_p2);

assign or_ln890_156_fu_38854_p2 = (xor_ln890_154_fu_38848_p2 | or_ln888_156_fu_38829_p2);

assign or_ln890_157_fu_39003_p2 = (xor_ln890_155_fu_38997_p2 | or_ln888_157_fu_38978_p2);

assign or_ln890_158_fu_39152_p2 = (xor_ln890_156_fu_39146_p2 | or_ln888_158_fu_39127_p2);

assign or_ln890_159_fu_34604_p2 = (xor_ln890_157_fu_34598_p2 | or_ln888_159_fu_34578_p2);

assign or_ln890_160_fu_39318_p2 = (xor_ln890_158_fu_39312_p2 | or_ln888_160_fu_39293_p2);

assign or_ln890_81_fu_19133_p2 = (xor_ln890_79_fu_19127_p2 | or_ln888_81_fu_19109_p2);

assign or_ln890_82_fu_19258_p2 = (xor_ln890_80_fu_19252_p2 | or_ln888_82_fu_19234_p2);

assign or_ln890_83_fu_19383_p2 = (xor_ln890_81_fu_19377_p2 | or_ln888_83_fu_19359_p2);

assign or_ln890_84_fu_19508_p2 = (xor_ln890_82_fu_19502_p2 | or_ln888_84_fu_19484_p2);

assign or_ln890_85_fu_19633_p2 = (xor_ln890_83_fu_19627_p2 | or_ln888_85_fu_19609_p2);

assign or_ln890_86_fu_19758_p2 = (xor_ln890_84_fu_19752_p2 | or_ln888_86_fu_19734_p2);

assign or_ln890_87_fu_19883_p2 = (xor_ln890_85_fu_19877_p2 | or_ln888_87_fu_19859_p2);

assign or_ln890_88_fu_20008_p2 = (xor_ln890_86_fu_20002_p2 | or_ln888_88_fu_19984_p2);

assign or_ln890_89_fu_20156_p2 = (xor_ln890_87_fu_20150_p2 | or_ln888_89_fu_20131_p2);

assign or_ln890_90_fu_20305_p2 = (xor_ln890_88_fu_20299_p2 | or_ln888_90_fu_20280_p2);

assign or_ln890_91_fu_20454_p2 = (xor_ln890_89_fu_20448_p2 | or_ln888_91_fu_20429_p2);

assign or_ln890_92_fu_20603_p2 = (xor_ln890_90_fu_20597_p2 | or_ln888_92_fu_20578_p2);

assign or_ln890_93_fu_20752_p2 = (xor_ln890_91_fu_20746_p2 | or_ln888_93_fu_20727_p2);

assign or_ln890_94_fu_18235_p2 = (xor_ln890_92_fu_18229_p2 | or_ln888_94_fu_18209_p2);

assign or_ln890_95_fu_20918_p2 = (xor_ln890_93_fu_20912_p2 | or_ln888_95_fu_20893_p2);

assign or_ln890_96_fu_21067_p2 = (xor_ln890_94_fu_21061_p2 | or_ln888_96_fu_21042_p2);

assign or_ln890_97_fu_21216_p2 = (xor_ln890_95_fu_21210_p2 | or_ln888_97_fu_21191_p2);

assign or_ln890_98_fu_21361_p2 = (xor_ln890_96_fu_21355_p2 | or_ln888_98_fu_21336_p2);

assign or_ln890_99_fu_21506_p2 = (xor_ln890_97_fu_21500_p2 | or_ln888_99_fu_21481_p2);

assign or_ln890_fu_19008_p2 = (xor_ln890_fu_19002_p2 | or_ln888_fu_18984_p2);

assign or_ln895_100_fu_21657_p2 = (xor_ln895_282_fu_21651_p2 | p_Result_464_fu_21586_p3);

assign or_ln895_101_fu_21782_p2 = (xor_ln895_284_fu_21776_p2 | p_Result_467_fu_21711_p3);

assign or_ln895_102_fu_21927_p2 = (xor_ln895_286_fu_21921_p2 | p_Result_470_fu_21856_p3);

assign or_ln895_103_fu_22056_p2 = (xor_ln895_288_fu_22050_p2 | p_Result_473_fu_21985_p3);

assign or_ln895_104_fu_22185_p2 = (xor_ln895_290_fu_22179_p2 | p_Result_476_fu_22114_p3);

assign or_ln895_105_fu_22314_p2 = (xor_ln895_292_fu_22308_p2 | p_Result_479_fu_22243_p3);

assign or_ln895_106_fu_22443_p2 = (xor_ln895_294_fu_22437_p2 | p_Result_482_fu_22372_p3);

assign or_ln895_107_fu_25605_p2 = (xor_ln895_296_fu_25599_p2 | p_Result_485_reg_42269);

assign or_ln895_108_fu_25730_p2 = (xor_ln895_298_fu_25724_p2 | p_Result_488_reg_42300);

assign or_ln895_109_fu_25855_p2 = (xor_ln895_300_fu_25849_p2 | p_Result_491_reg_42331);

assign or_ln895_110_fu_25980_p2 = (xor_ln895_302_fu_25974_p2 | p_Result_494_reg_42362);

assign or_ln895_111_fu_26105_p2 = (xor_ln895_304_fu_26099_p2 | p_Result_497_reg_42393);

assign or_ln895_112_fu_26230_p2 = (xor_ln895_306_fu_26224_p2 | p_Result_500_reg_42424);

assign or_ln895_113_fu_23041_p2 = (xor_ln895_308_fu_23035_p2 | p_Result_503_fu_22957_p3);

assign or_ln895_114_fu_26372_p2 = (xor_ln895_310_fu_26366_p2 | p_Result_506_reg_42470);

assign or_ln895_115_fu_26497_p2 = (xor_ln895_312_fu_26491_p2 | p_Result_509_reg_42501);

assign or_ln895_116_fu_26641_p2 = (xor_ln895_314_fu_26635_p2 | p_Result_512_fu_26570_p3);

assign or_ln895_117_fu_26790_p2 = (xor_ln895_316_fu_26784_p2 | p_Result_515_fu_26719_p3);

assign or_ln895_118_fu_26939_p2 = (xor_ln895_318_fu_26933_p2 | p_Result_518_fu_26868_p3);

assign or_ln895_119_fu_27088_p2 = (xor_ln895_320_fu_27082_p2 | p_Result_521_fu_27017_p3);

assign or_ln895_120_fu_27237_p2 = (xor_ln895_322_fu_27231_p2 | p_Result_524_fu_27166_p3);

assign or_ln895_121_fu_27386_p2 = (xor_ln895_324_fu_27380_p2 | p_Result_527_fu_27315_p3);

assign or_ln895_122_fu_27535_p2 = (xor_ln895_326_fu_27529_p2 | p_Result_530_fu_27464_p3);

assign or_ln895_123_fu_27684_p2 = (xor_ln895_328_fu_27678_p2 | p_Result_533_fu_27613_p3);

assign or_ln895_124_fu_27833_p2 = (xor_ln895_330_fu_27827_p2 | p_Result_536_fu_27762_p3);

assign or_ln895_125_fu_28069_p2 = (xor_ln895_332_fu_28063_p2 | p_Result_539_fu_27985_p3);

assign or_ln895_126_fu_31403_p2 = (xor_ln895_334_fu_31397_p2 | p_Result_542_reg_42862);

assign or_ln895_127_fu_31528_p2 = (xor_ln895_336_fu_31522_p2 | p_Result_545_reg_42893);

assign or_ln895_128_fu_31653_p2 = (xor_ln895_338_fu_31647_p2 | p_Result_548_reg_42924);

assign or_ln895_129_fu_31778_p2 = (xor_ln895_340_fu_31772_p2 | p_Result_551_reg_42955);

assign or_ln895_130_fu_31903_p2 = (xor_ln895_342_fu_31897_p2 | p_Result_554_reg_42986);

assign or_ln895_131_fu_32028_p2 = (xor_ln895_344_fu_32022_p2 | p_Result_557_reg_43017);

assign or_ln895_132_fu_32153_p2 = (xor_ln895_346_fu_32147_p2 | p_Result_560_reg_43048);

assign or_ln895_133_fu_32278_p2 = (xor_ln895_348_fu_32272_p2 | p_Result_563_reg_43079);

assign or_ln895_134_fu_32426_p2 = (xor_ln895_350_fu_32420_p2 | p_Result_566_fu_32355_p3);

assign or_ln895_135_fu_32575_p2 = (xor_ln895_352_fu_32569_p2 | p_Result_569_fu_32504_p3);

assign or_ln895_136_fu_32724_p2 = (xor_ln895_354_fu_32718_p2 | p_Result_572_fu_32653_p3);

assign or_ln895_137_fu_32873_p2 = (xor_ln895_356_fu_32867_p2 | p_Result_575_fu_32802_p3);

assign or_ln895_138_fu_33022_p2 = (xor_ln895_358_fu_33016_p2 | p_Result_578_fu_32951_p3);

assign or_ln895_139_fu_33171_p2 = (xor_ln895_360_fu_33165_p2 | p_Result_581_fu_33100_p3);

assign or_ln895_140_fu_33320_p2 = (xor_ln895_362_fu_33314_p2 | p_Result_584_fu_33249_p3);

assign or_ln895_141_fu_33469_p2 = (xor_ln895_364_fu_33463_p2 | p_Result_587_fu_33398_p3);

assign or_ln895_142_fu_29136_p2 = (xor_ln895_366_fu_29130_p2 | p_Result_590_fu_29052_p3);

assign or_ln895_143_fu_37137_p2 = (xor_ln895_368_fu_37131_p2 | p_Result_593_reg_43537);

assign or_ln895_144_fu_37261_p2 = (xor_ln895_370_fu_37255_p2 | p_Result_596_reg_43568);

assign or_ln895_145_fu_37386_p2 = (xor_ln895_372_fu_37380_p2 | p_Result_599_reg_43599);

assign or_ln895_146_fu_37511_p2 = (xor_ln895_374_fu_37505_p2 | p_Result_602_reg_43630);

assign or_ln895_147_fu_37636_p2 = (xor_ln895_376_fu_37630_p2 | p_Result_605_reg_43661);

assign or_ln895_148_fu_37761_p2 = (xor_ln895_378_fu_37755_p2 | p_Result_608_reg_43692);

assign or_ln895_149_fu_37886_p2 = (xor_ln895_380_fu_37880_p2 | p_Result_611_reg_43723);

assign or_ln895_150_fu_38011_p2 = (xor_ln895_382_fu_38005_p2 | p_Result_614_reg_43754);

assign or_ln895_151_fu_38136_p2 = (xor_ln895_384_fu_38130_p2 | p_Result_617_reg_43785);

assign or_ln895_152_fu_38280_p2 = (xor_ln895_386_fu_38274_p2 | p_Result_620_fu_38209_p3);

assign or_ln895_153_fu_38429_p2 = (xor_ln895_388_fu_38423_p2 | p_Result_623_fu_38358_p3);

assign or_ln895_154_fu_38578_p2 = (xor_ln895_390_fu_38572_p2 | p_Result_626_fu_38507_p3);

assign or_ln895_155_fu_38727_p2 = (xor_ln895_392_fu_38721_p2 | p_Result_629_fu_38656_p3);

assign or_ln895_156_fu_38876_p2 = (xor_ln895_394_fu_38870_p2 | p_Result_632_fu_38805_p3);

assign or_ln895_157_fu_39025_p2 = (xor_ln895_396_fu_39019_p2 | p_Result_635_fu_38954_p3);

assign or_ln895_158_fu_39174_p2 = (xor_ln895_398_fu_39168_p2 | p_Result_638_fu_39103_p3);

assign or_ln895_159_fu_34628_p2 = (xor_ln895_400_fu_34622_p2 | p_Result_641_fu_34544_p3);

assign or_ln895_160_fu_39340_p2 = (xor_ln895_402_fu_39334_p2 | p_Result_644_fu_39269_p3);

assign or_ln895_81_fu_19155_p2 = (xor_ln895_244_fu_19149_p2 | p_Result_407_reg_41381);

assign or_ln895_82_fu_19280_p2 = (xor_ln895_246_fu_19274_p2 | p_Result_410_reg_41412);

assign or_ln895_83_fu_19405_p2 = (xor_ln895_248_fu_19399_p2 | p_Result_413_reg_41443);

assign or_ln895_84_fu_19530_p2 = (xor_ln895_250_fu_19524_p2 | p_Result_416_reg_41474);

assign or_ln895_85_fu_19655_p2 = (xor_ln895_252_fu_19649_p2 | p_Result_419_reg_41505);

assign or_ln895_86_fu_19780_p2 = (xor_ln895_254_fu_19774_p2 | p_Result_422_reg_41536);

assign or_ln895_87_fu_19905_p2 = (xor_ln895_256_fu_19899_p2 | p_Result_425_reg_41567);

assign or_ln895_88_fu_20030_p2 = (xor_ln895_258_fu_20024_p2 | p_Result_428_reg_41598);

assign or_ln895_89_fu_20178_p2 = (xor_ln895_260_fu_20172_p2 | p_Result_431_fu_20107_p3);

assign or_ln895_90_fu_20327_p2 = (xor_ln895_262_fu_20321_p2 | p_Result_434_fu_20256_p3);

assign or_ln895_91_fu_20476_p2 = (xor_ln895_264_fu_20470_p2 | p_Result_437_fu_20405_p3);

assign or_ln895_92_fu_20625_p2 = (xor_ln895_266_fu_20619_p2 | p_Result_440_fu_20554_p3);

assign or_ln895_93_fu_20774_p2 = (xor_ln895_268_fu_20768_p2 | p_Result_443_fu_20703_p3);

assign or_ln895_94_fu_18259_p2 = (xor_ln895_270_fu_18253_p2 | p_Result_446_fu_18175_p3);

assign or_ln895_95_fu_20940_p2 = (xor_ln895_272_fu_20934_p2 | p_Result_449_fu_20869_p3);

assign or_ln895_96_fu_21089_p2 = (xor_ln895_274_fu_21083_p2 | p_Result_452_fu_21018_p3);

assign or_ln895_97_fu_21238_p2 = (xor_ln895_276_fu_21232_p2 | p_Result_455_fu_21167_p3);

assign or_ln895_98_fu_21383_p2 = (xor_ln895_278_fu_21377_p2 | p_Result_458_fu_21312_p3);

assign or_ln895_99_fu_21528_p2 = (xor_ln895_280_fu_21522_p2 | p_Result_461_fu_21457_p3);

assign or_ln895_fu_19030_p2 = (xor_ln895_fu_19024_p2 | p_Result_404_reg_41350);

assign or_ln896_100_fu_21680_p2 = (xor_ln896_283_fu_21674_p2 | xor_ln896_282_fu_21594_p2);

assign or_ln896_101_fu_21805_p2 = (xor_ln896_285_fu_21799_p2 | xor_ln896_284_fu_21719_p2);

assign or_ln896_102_fu_21950_p2 = (xor_ln896_287_fu_21944_p2 | xor_ln896_286_fu_21864_p2);

assign or_ln896_103_fu_22079_p2 = (xor_ln896_289_fu_22073_p2 | xor_ln896_288_fu_21993_p2);

assign or_ln896_104_fu_22208_p2 = (xor_ln896_291_fu_22202_p2 | xor_ln896_290_fu_22122_p2);

assign or_ln896_105_fu_22337_p2 = (xor_ln896_293_fu_22331_p2 | xor_ln896_292_fu_22251_p2);

assign or_ln896_106_fu_22466_p2 = (xor_ln896_295_fu_22460_p2 | xor_ln896_294_fu_22380_p2);

assign or_ln896_107_fu_25627_p2 = (xor_ln896_297_fu_25621_p2 | xor_ln896_296_fu_25544_p2);

assign or_ln896_108_fu_25752_p2 = (xor_ln896_299_fu_25746_p2 | xor_ln896_298_fu_25669_p2);

assign or_ln896_109_fu_25877_p2 = (xor_ln896_301_fu_25871_p2 | xor_ln896_300_fu_25794_p2);

assign or_ln896_110_fu_26002_p2 = (xor_ln896_303_fu_25996_p2 | xor_ln896_302_fu_25919_p2);

assign or_ln896_111_fu_26127_p2 = (xor_ln896_305_fu_26121_p2 | xor_ln896_304_fu_26044_p2);

assign or_ln896_112_fu_26252_p2 = (xor_ln896_307_fu_26246_p2 | xor_ln896_306_fu_26169_p2);

assign or_ln896_113_fu_23065_p2 = (xor_ln896_309_fu_23059_p2 | xor_ln896_308_fu_22965_p2);

assign or_ln896_114_fu_26394_p2 = (xor_ln896_311_fu_26388_p2 | xor_ln896_310_fu_26311_p2);

assign or_ln896_115_fu_26519_p2 = (xor_ln896_313_fu_26513_p2 | xor_ln896_312_fu_26436_p2);

assign or_ln896_116_fu_26664_p2 = (xor_ln896_315_fu_26658_p2 | xor_ln896_314_fu_26578_p2);

assign or_ln896_117_fu_26813_p2 = (xor_ln896_317_fu_26807_p2 | xor_ln896_316_fu_26727_p2);

assign or_ln896_118_fu_26962_p2 = (xor_ln896_319_fu_26956_p2 | xor_ln896_318_fu_26876_p2);

assign or_ln896_119_fu_27111_p2 = (xor_ln896_321_fu_27105_p2 | xor_ln896_320_fu_27025_p2);

assign or_ln896_120_fu_27260_p2 = (xor_ln896_323_fu_27254_p2 | xor_ln896_322_fu_27174_p2);

assign or_ln896_121_fu_27409_p2 = (xor_ln896_325_fu_27403_p2 | xor_ln896_324_fu_27323_p2);

assign or_ln896_122_fu_27558_p2 = (xor_ln896_327_fu_27552_p2 | xor_ln896_326_fu_27472_p2);

assign or_ln896_123_fu_27707_p2 = (xor_ln896_329_fu_27701_p2 | xor_ln896_328_fu_27621_p2);

assign or_ln896_124_fu_27856_p2 = (xor_ln896_331_fu_27850_p2 | xor_ln896_330_fu_27770_p2);

assign or_ln896_125_fu_28093_p2 = (xor_ln896_333_fu_28087_p2 | xor_ln896_332_fu_27993_p2);

assign or_ln896_126_fu_31425_p2 = (xor_ln896_335_fu_31419_p2 | xor_ln896_334_fu_31342_p2);

assign or_ln896_127_fu_31550_p2 = (xor_ln896_337_fu_31544_p2 | xor_ln896_336_fu_31467_p2);

assign or_ln896_128_fu_31675_p2 = (xor_ln896_339_fu_31669_p2 | xor_ln896_338_fu_31592_p2);

assign or_ln896_129_fu_31800_p2 = (xor_ln896_341_fu_31794_p2 | xor_ln896_340_fu_31717_p2);

assign or_ln896_130_fu_31925_p2 = (xor_ln896_343_fu_31919_p2 | xor_ln896_342_fu_31842_p2);

assign or_ln896_131_fu_32050_p2 = (xor_ln896_345_fu_32044_p2 | xor_ln896_344_fu_31967_p2);

assign or_ln896_132_fu_32175_p2 = (xor_ln896_347_fu_32169_p2 | xor_ln896_346_fu_32092_p2);

assign or_ln896_133_fu_32300_p2 = (xor_ln896_349_fu_32294_p2 | xor_ln896_348_fu_32217_p2);

assign or_ln896_134_fu_32449_p2 = (xor_ln896_351_fu_32443_p2 | xor_ln896_350_fu_32363_p2);

assign or_ln896_135_fu_32598_p2 = (xor_ln896_353_fu_32592_p2 | xor_ln896_352_fu_32512_p2);

assign or_ln896_136_fu_32747_p2 = (xor_ln896_355_fu_32741_p2 | xor_ln896_354_fu_32661_p2);

assign or_ln896_137_fu_32896_p2 = (xor_ln896_357_fu_32890_p2 | xor_ln896_356_fu_32810_p2);

assign or_ln896_138_fu_33045_p2 = (xor_ln896_359_fu_33039_p2 | xor_ln896_358_fu_32959_p2);

assign or_ln896_139_fu_33194_p2 = (xor_ln896_361_fu_33188_p2 | xor_ln896_360_fu_33108_p2);

assign or_ln896_140_fu_33343_p2 = (xor_ln896_363_fu_33337_p2 | xor_ln896_362_fu_33257_p2);

assign or_ln896_141_fu_33492_p2 = (xor_ln896_365_fu_33486_p2 | xor_ln896_364_fu_33406_p2);

assign or_ln896_142_fu_29160_p2 = (xor_ln896_367_fu_29154_p2 | xor_ln896_366_fu_29060_p2);

assign or_ln896_143_fu_37159_p2 = (xor_ln896_369_fu_37153_p2 | xor_ln896_368_fu_37076_p2);

assign or_ln896_144_fu_37283_p2 = (xor_ln896_371_fu_37277_p2 | xor_ln896_370_fu_37200_p2);

assign or_ln896_145_fu_37408_p2 = (xor_ln896_373_fu_37402_p2 | xor_ln896_372_fu_37325_p2);

assign or_ln896_146_fu_37533_p2 = (xor_ln896_375_fu_37527_p2 | xor_ln896_374_fu_37450_p2);

assign or_ln896_147_fu_37658_p2 = (xor_ln896_377_fu_37652_p2 | xor_ln896_376_fu_37575_p2);

assign or_ln896_148_fu_37783_p2 = (xor_ln896_379_fu_37777_p2 | xor_ln896_378_fu_37700_p2);

assign or_ln896_149_fu_37908_p2 = (xor_ln896_381_fu_37902_p2 | xor_ln896_380_fu_37825_p2);

assign or_ln896_150_fu_38033_p2 = (xor_ln896_383_fu_38027_p2 | xor_ln896_382_fu_37950_p2);

assign or_ln896_151_fu_38158_p2 = (xor_ln896_385_fu_38152_p2 | xor_ln896_384_fu_38075_p2);

assign or_ln896_152_fu_38303_p2 = (xor_ln896_387_fu_38297_p2 | xor_ln896_386_fu_38217_p2);

assign or_ln896_153_fu_38452_p2 = (xor_ln896_389_fu_38446_p2 | xor_ln896_388_fu_38366_p2);

assign or_ln896_154_fu_38601_p2 = (xor_ln896_391_fu_38595_p2 | xor_ln896_390_fu_38515_p2);

assign or_ln896_155_fu_38750_p2 = (xor_ln896_393_fu_38744_p2 | xor_ln896_392_fu_38664_p2);

assign or_ln896_156_fu_38899_p2 = (xor_ln896_395_fu_38893_p2 | xor_ln896_394_fu_38813_p2);

assign or_ln896_157_fu_39048_p2 = (xor_ln896_397_fu_39042_p2 | xor_ln896_396_fu_38962_p2);

assign or_ln896_158_fu_39197_p2 = (xor_ln896_399_fu_39191_p2 | xor_ln896_398_fu_39111_p2);

assign or_ln896_159_fu_34652_p2 = (xor_ln896_401_fu_34646_p2 | xor_ln896_400_fu_34552_p2);

assign or_ln896_160_fu_39363_p2 = (xor_ln896_403_fu_39357_p2 | xor_ln896_402_fu_39277_p2);

assign or_ln896_81_fu_19177_p2 = (xor_ln896_245_fu_19171_p2 | xor_ln896_244_fu_19094_p2);

assign or_ln896_82_fu_19302_p2 = (xor_ln896_247_fu_19296_p2 | xor_ln896_246_fu_19219_p2);

assign or_ln896_83_fu_19427_p2 = (xor_ln896_249_fu_19421_p2 | xor_ln896_248_fu_19344_p2);

assign or_ln896_84_fu_19552_p2 = (xor_ln896_251_fu_19546_p2 | xor_ln896_250_fu_19469_p2);

assign or_ln896_85_fu_19677_p2 = (xor_ln896_253_fu_19671_p2 | xor_ln896_252_fu_19594_p2);

assign or_ln896_86_fu_19802_p2 = (xor_ln896_255_fu_19796_p2 | xor_ln896_254_fu_19719_p2);

assign or_ln896_87_fu_19927_p2 = (xor_ln896_257_fu_19921_p2 | xor_ln896_256_fu_19844_p2);

assign or_ln896_88_fu_20052_p2 = (xor_ln896_259_fu_20046_p2 | xor_ln896_258_fu_19969_p2);

assign or_ln896_89_fu_20201_p2 = (xor_ln896_261_fu_20195_p2 | xor_ln896_260_fu_20115_p2);

assign or_ln896_90_fu_20350_p2 = (xor_ln896_263_fu_20344_p2 | xor_ln896_262_fu_20264_p2);

assign or_ln896_91_fu_20499_p2 = (xor_ln896_265_fu_20493_p2 | xor_ln896_264_fu_20413_p2);

assign or_ln896_92_fu_20648_p2 = (xor_ln896_267_fu_20642_p2 | xor_ln896_266_fu_20562_p2);

assign or_ln896_93_fu_20797_p2 = (xor_ln896_269_fu_20791_p2 | xor_ln896_268_fu_20711_p2);

assign or_ln896_94_fu_18283_p2 = (xor_ln896_271_fu_18277_p2 | xor_ln896_270_fu_18183_p2);

assign or_ln896_95_fu_20963_p2 = (xor_ln896_273_fu_20957_p2 | xor_ln896_272_fu_20877_p2);

assign or_ln896_96_fu_21112_p2 = (xor_ln896_275_fu_21106_p2 | xor_ln896_274_fu_21026_p2);

assign or_ln896_97_fu_21261_p2 = (xor_ln896_277_fu_21255_p2 | xor_ln896_276_fu_21175_p2);

assign or_ln896_98_fu_21406_p2 = (xor_ln896_279_fu_21400_p2 | xor_ln896_278_fu_21320_p2);

assign or_ln896_99_fu_21551_p2 = (xor_ln896_281_fu_21545_p2 | xor_ln896_280_fu_21465_p2);

assign or_ln896_fu_19052_p2 = (xor_ln896_fu_18969_p2 | xor_ln896_243_fu_19046_p2);

assign overflow_162_fu_19165_p2 = (xor_ln895_245_fu_19160_p2 & or_ln895_81_fu_19155_p2);

assign overflow_163_fu_19290_p2 = (xor_ln895_247_fu_19285_p2 & or_ln895_82_fu_19280_p2);

assign overflow_164_fu_19415_p2 = (xor_ln895_249_fu_19410_p2 & or_ln895_83_fu_19405_p2);

assign overflow_165_fu_19540_p2 = (xor_ln895_251_fu_19535_p2 & or_ln895_84_fu_19530_p2);

assign overflow_166_fu_19665_p2 = (xor_ln895_253_fu_19660_p2 & or_ln895_85_fu_19655_p2);

assign overflow_167_fu_19790_p2 = (xor_ln895_255_fu_19785_p2 & or_ln895_86_fu_19780_p2);

assign overflow_168_fu_19915_p2 = (xor_ln895_257_fu_19910_p2 & or_ln895_87_fu_19905_p2);

assign overflow_169_fu_20040_p2 = (xor_ln895_259_fu_20035_p2 & or_ln895_88_fu_20030_p2);

assign overflow_170_fu_20189_p2 = (xor_ln895_261_fu_20184_p2 & or_ln895_89_fu_20178_p2);

assign overflow_171_fu_20338_p2 = (xor_ln895_263_fu_20333_p2 & or_ln895_90_fu_20327_p2);

assign overflow_172_fu_20487_p2 = (xor_ln895_265_fu_20482_p2 & or_ln895_91_fu_20476_p2);

assign overflow_173_fu_20636_p2 = (xor_ln895_267_fu_20631_p2 & or_ln895_92_fu_20625_p2);

assign overflow_174_fu_20785_p2 = (xor_ln895_269_fu_20780_p2 & or_ln895_93_fu_20774_p2);

assign overflow_175_fu_18271_p2 = (xor_ln895_271_fu_18265_p2 & or_ln895_94_fu_18259_p2);

assign overflow_176_fu_20951_p2 = (xor_ln895_273_fu_20946_p2 & or_ln895_95_fu_20940_p2);

assign overflow_177_fu_21100_p2 = (xor_ln895_275_fu_21095_p2 & or_ln895_96_fu_21089_p2);

assign overflow_178_fu_21249_p2 = (xor_ln895_277_fu_21244_p2 & or_ln895_97_fu_21238_p2);

assign overflow_179_fu_21394_p2 = (xor_ln895_279_fu_21389_p2 & or_ln895_98_fu_21383_p2);

assign overflow_180_fu_21539_p2 = (xor_ln895_281_fu_21534_p2 & or_ln895_99_fu_21528_p2);

assign overflow_181_fu_21668_p2 = (xor_ln895_283_fu_21663_p2 & or_ln895_100_fu_21657_p2);

assign overflow_182_fu_21793_p2 = (xor_ln895_285_fu_21788_p2 & or_ln895_101_fu_21782_p2);

assign overflow_183_fu_21938_p2 = (xor_ln895_287_fu_21933_p2 & or_ln895_102_fu_21927_p2);

assign overflow_184_fu_22067_p2 = (xor_ln895_289_fu_22062_p2 & or_ln895_103_fu_22056_p2);

assign overflow_185_fu_22196_p2 = (xor_ln895_291_fu_22191_p2 & or_ln895_104_fu_22185_p2);

assign overflow_186_fu_22325_p2 = (xor_ln895_293_fu_22320_p2 & or_ln895_105_fu_22314_p2);

assign overflow_187_fu_22454_p2 = (xor_ln895_295_fu_22449_p2 & or_ln895_106_fu_22443_p2);

assign overflow_188_fu_25615_p2 = (xor_ln895_297_fu_25610_p2 & or_ln895_107_fu_25605_p2);

assign overflow_189_fu_25740_p2 = (xor_ln895_299_fu_25735_p2 & or_ln895_108_fu_25730_p2);

assign overflow_190_fu_25865_p2 = (xor_ln895_301_fu_25860_p2 & or_ln895_109_fu_25855_p2);

assign overflow_191_fu_25990_p2 = (xor_ln895_303_fu_25985_p2 & or_ln895_110_fu_25980_p2);

assign overflow_192_fu_26115_p2 = (xor_ln895_305_fu_26110_p2 & or_ln895_111_fu_26105_p2);

assign overflow_193_fu_26240_p2 = (xor_ln895_307_fu_26235_p2 & or_ln895_112_fu_26230_p2);

assign overflow_194_fu_23053_p2 = (xor_ln895_309_fu_23047_p2 & or_ln895_113_fu_23041_p2);

assign overflow_195_fu_26382_p2 = (xor_ln895_311_fu_26377_p2 & or_ln895_114_fu_26372_p2);

assign overflow_196_fu_26507_p2 = (xor_ln895_313_fu_26502_p2 & or_ln895_115_fu_26497_p2);

assign overflow_197_fu_26652_p2 = (xor_ln895_315_fu_26647_p2 & or_ln895_116_fu_26641_p2);

assign overflow_198_fu_26801_p2 = (xor_ln895_317_fu_26796_p2 & or_ln895_117_fu_26790_p2);

assign overflow_199_fu_26950_p2 = (xor_ln895_319_fu_26945_p2 & or_ln895_118_fu_26939_p2);

assign overflow_200_fu_27099_p2 = (xor_ln895_321_fu_27094_p2 & or_ln895_119_fu_27088_p2);

assign overflow_201_fu_27248_p2 = (xor_ln895_323_fu_27243_p2 & or_ln895_120_fu_27237_p2);

assign overflow_202_fu_27397_p2 = (xor_ln895_325_fu_27392_p2 & or_ln895_121_fu_27386_p2);

assign overflow_203_fu_27546_p2 = (xor_ln895_327_fu_27541_p2 & or_ln895_122_fu_27535_p2);

assign overflow_204_fu_27695_p2 = (xor_ln895_329_fu_27690_p2 & or_ln895_123_fu_27684_p2);

assign overflow_205_fu_27844_p2 = (xor_ln895_331_fu_27839_p2 & or_ln895_124_fu_27833_p2);

assign overflow_206_fu_28081_p2 = (xor_ln895_333_fu_28075_p2 & or_ln895_125_fu_28069_p2);

assign overflow_207_fu_31413_p2 = (xor_ln895_335_fu_31408_p2 & or_ln895_126_fu_31403_p2);

assign overflow_208_fu_31538_p2 = (xor_ln895_337_fu_31533_p2 & or_ln895_127_fu_31528_p2);

assign overflow_209_fu_31663_p2 = (xor_ln895_339_fu_31658_p2 & or_ln895_128_fu_31653_p2);

assign overflow_210_fu_31788_p2 = (xor_ln895_341_fu_31783_p2 & or_ln895_129_fu_31778_p2);

assign overflow_211_fu_31913_p2 = (xor_ln895_343_fu_31908_p2 & or_ln895_130_fu_31903_p2);

assign overflow_212_fu_32038_p2 = (xor_ln895_345_fu_32033_p2 & or_ln895_131_fu_32028_p2);

assign overflow_213_fu_32163_p2 = (xor_ln895_347_fu_32158_p2 & or_ln895_132_fu_32153_p2);

assign overflow_214_fu_32288_p2 = (xor_ln895_349_fu_32283_p2 & or_ln895_133_fu_32278_p2);

assign overflow_215_fu_32437_p2 = (xor_ln895_351_fu_32432_p2 & or_ln895_134_fu_32426_p2);

assign overflow_216_fu_32586_p2 = (xor_ln895_353_fu_32581_p2 & or_ln895_135_fu_32575_p2);

assign overflow_217_fu_32735_p2 = (xor_ln895_355_fu_32730_p2 & or_ln895_136_fu_32724_p2);

assign overflow_218_fu_32884_p2 = (xor_ln895_357_fu_32879_p2 & or_ln895_137_fu_32873_p2);

assign overflow_219_fu_33033_p2 = (xor_ln895_359_fu_33028_p2 & or_ln895_138_fu_33022_p2);

assign overflow_220_fu_33182_p2 = (xor_ln895_361_fu_33177_p2 & or_ln895_139_fu_33171_p2);

assign overflow_221_fu_33331_p2 = (xor_ln895_363_fu_33326_p2 & or_ln895_140_fu_33320_p2);

assign overflow_222_fu_33480_p2 = (xor_ln895_365_fu_33475_p2 & or_ln895_141_fu_33469_p2);

assign overflow_223_fu_29148_p2 = (xor_ln895_367_fu_29142_p2 & or_ln895_142_fu_29136_p2);

assign overflow_224_fu_37147_p2 = (xor_ln895_369_fu_37142_p2 & or_ln895_143_fu_37137_p2);

assign overflow_225_fu_37271_p2 = (xor_ln895_371_fu_37266_p2 & or_ln895_144_fu_37261_p2);

assign overflow_226_fu_37396_p2 = (xor_ln895_373_fu_37391_p2 & or_ln895_145_fu_37386_p2);

assign overflow_227_fu_37521_p2 = (xor_ln895_375_fu_37516_p2 & or_ln895_146_fu_37511_p2);

assign overflow_228_fu_37646_p2 = (xor_ln895_377_fu_37641_p2 & or_ln895_147_fu_37636_p2);

assign overflow_229_fu_37771_p2 = (xor_ln895_379_fu_37766_p2 & or_ln895_148_fu_37761_p2);

assign overflow_230_fu_37896_p2 = (xor_ln895_381_fu_37891_p2 & or_ln895_149_fu_37886_p2);

assign overflow_231_fu_38021_p2 = (xor_ln895_383_fu_38016_p2 & or_ln895_150_fu_38011_p2);

assign overflow_232_fu_38146_p2 = (xor_ln895_385_fu_38141_p2 & or_ln895_151_fu_38136_p2);

assign overflow_233_fu_38291_p2 = (xor_ln895_387_fu_38286_p2 & or_ln895_152_fu_38280_p2);

assign overflow_234_fu_38440_p2 = (xor_ln895_389_fu_38435_p2 & or_ln895_153_fu_38429_p2);

assign overflow_235_fu_38589_p2 = (xor_ln895_391_fu_38584_p2 & or_ln895_154_fu_38578_p2);

assign overflow_236_fu_38738_p2 = (xor_ln895_393_fu_38733_p2 & or_ln895_155_fu_38727_p2);

assign overflow_237_fu_38887_p2 = (xor_ln895_395_fu_38882_p2 & or_ln895_156_fu_38876_p2);

assign overflow_238_fu_39036_p2 = (xor_ln895_397_fu_39031_p2 & or_ln895_157_fu_39025_p2);

assign overflow_239_fu_39185_p2 = (xor_ln895_399_fu_39180_p2 & or_ln895_158_fu_39174_p2);

assign overflow_240_fu_34640_p2 = (xor_ln895_401_fu_34634_p2 & or_ln895_159_fu_34628_p2);

assign overflow_241_fu_39351_p2 = (xor_ln895_403_fu_39346_p2 & or_ln895_160_fu_39340_p2);

assign overflow_242_fu_23660_p2 = (xor_ln895_404_fu_23654_p2 & p_Result_646_fu_23646_p3);

assign overflow_243_fu_23758_p2 = (xor_ln895_405_fu_23752_p2 & p_Result_648_fu_23744_p3);

assign overflow_244_fu_23856_p2 = (xor_ln895_406_fu_23850_p2 & p_Result_650_fu_23842_p3);

assign overflow_245_fu_23954_p2 = (xor_ln895_407_fu_23948_p2 & p_Result_652_fu_23940_p3);

assign overflow_246_fu_24052_p2 = (xor_ln895_408_fu_24046_p2 & p_Result_654_fu_24038_p3);

assign overflow_247_fu_24150_p2 = (xor_ln895_409_fu_24144_p2 & p_Result_656_fu_24136_p3);

assign overflow_248_fu_24248_p2 = (xor_ln895_410_fu_24242_p2 & p_Result_658_fu_24234_p3);

assign overflow_249_fu_24346_p2 = (xor_ln895_411_fu_24340_p2 & p_Result_660_fu_24332_p3);

assign overflow_250_fu_24444_p2 = (xor_ln895_412_fu_24438_p2 & p_Result_662_fu_24430_p3);

assign overflow_251_fu_24546_p2 = (xor_ln895_413_fu_24540_p2 & p_Result_664_fu_24532_p3);

assign overflow_252_fu_24648_p2 = (xor_ln895_414_fu_24642_p2 & p_Result_666_fu_24634_p3);

assign overflow_253_fu_24750_p2 = (xor_ln895_415_fu_24744_p2 & p_Result_668_fu_24736_p3);

assign overflow_254_fu_24852_p2 = (xor_ln895_416_fu_24846_p2 & p_Result_670_fu_24838_p3);

assign overflow_255_fu_24954_p2 = (xor_ln895_417_fu_24948_p2 & p_Result_672_fu_24940_p3);

assign overflow_256_fu_25056_p2 = (xor_ln895_418_fu_25050_p2 & p_Result_674_fu_25042_p3);

assign overflow_257_fu_25158_p2 = (xor_ln895_419_fu_25152_p2 & p_Result_676_fu_25144_p3);

assign overflow_258_fu_25260_p2 = (xor_ln895_420_fu_25254_p2 & p_Result_678_fu_25246_p3);

assign overflow_259_fu_25362_p2 = (xor_ln895_421_fu_25356_p2 & p_Result_680_fu_25348_p3);

assign overflow_260_fu_29222_p2 = (xor_ln895_422_fu_29216_p2 & p_Result_682_fu_29208_p3);

assign overflow_261_fu_29322_p2 = (xor_ln895_423_fu_29316_p2 & p_Result_684_fu_29308_p3);

assign overflow_262_fu_29422_p2 = (xor_ln895_424_fu_29416_p2 & p_Result_686_fu_29408_p3);

assign overflow_263_fu_29520_p2 = (xor_ln895_425_fu_29514_p2 & p_Result_688_fu_29506_p3);

assign overflow_264_fu_29620_p2 = (xor_ln895_426_fu_29614_p2 & p_Result_690_fu_29606_p3);

assign overflow_265_fu_29720_p2 = (xor_ln895_427_fu_29714_p2 & p_Result_692_fu_29706_p3);

assign overflow_266_fu_29820_p2 = (xor_ln895_428_fu_29814_p2 & p_Result_694_fu_29806_p3);

assign overflow_267_fu_29920_p2 = (xor_ln895_429_fu_29914_p2 & p_Result_696_fu_29906_p3);

assign overflow_268_fu_30020_p2 = (xor_ln895_430_fu_30014_p2 & p_Result_698_fu_30006_p3);

assign overflow_269_fu_30122_p2 = (xor_ln895_431_fu_30116_p2 & p_Result_700_fu_30108_p3);

assign overflow_270_fu_30224_p2 = (xor_ln895_432_fu_30218_p2 & p_Result_702_fu_30210_p3);

assign overflow_271_fu_30326_p2 = (xor_ln895_433_fu_30320_p2 & p_Result_704_fu_30312_p3);

assign overflow_272_fu_30428_p2 = (xor_ln895_434_fu_30422_p2 & p_Result_706_fu_30414_p3);

assign overflow_273_fu_30530_p2 = (xor_ln895_435_fu_30524_p2 & p_Result_708_fu_30516_p3);

assign overflow_274_fu_30632_p2 = (xor_ln895_436_fu_30626_p2 & p_Result_710_fu_30618_p3);

assign overflow_275_fu_30734_p2 = (xor_ln895_437_fu_30728_p2 & p_Result_712_fu_30720_p3);

assign overflow_276_fu_30836_p2 = (xor_ln895_438_fu_30830_p2 & p_Result_714_fu_30822_p3);

assign overflow_277_fu_30938_p2 = (xor_ln895_439_fu_30932_p2 & p_Result_716_fu_30924_p3);

assign overflow_278_fu_34723_p2 = (xor_ln895_440_fu_34718_p2 & p_Result_718_reg_43353);

assign overflow_279_fu_34781_p2 = (xor_ln895_441_fu_34776_p2 & p_Result_720_reg_43373);

assign overflow_280_fu_34839_p2 = (xor_ln895_442_fu_34834_p2 & p_Result_722_reg_43393);

assign overflow_281_fu_34897_p2 = (xor_ln895_443_fu_34892_p2 & p_Result_724_reg_43413);

assign overflow_282_fu_34955_p2 = (xor_ln895_444_fu_34950_p2 & p_Result_726_reg_43433);

assign overflow_283_fu_35013_p2 = (xor_ln895_445_fu_35008_p2 & p_Result_728_reg_43453);

assign overflow_284_fu_35071_p2 = (xor_ln895_446_fu_35066_p2 & p_Result_730_reg_43473);

assign overflow_285_fu_35129_p2 = (xor_ln895_447_fu_35124_p2 & p_Result_732_reg_43493);

assign overflow_286_fu_35187_p2 = (xor_ln895_448_fu_35182_p2 & p_Result_734_reg_43513);

assign overflow_287_fu_35282_p2 = (xor_ln895_449_fu_35276_p2 & p_Result_736_fu_35268_p3);

assign overflow_288_fu_35384_p2 = (xor_ln895_450_fu_35378_p2 & p_Result_738_fu_35370_p3);

assign overflow_289_fu_35486_p2 = (xor_ln895_451_fu_35480_p2 & p_Result_740_fu_35472_p3);

assign overflow_290_fu_35588_p2 = (xor_ln895_452_fu_35582_p2 & p_Result_742_fu_35574_p3);

assign overflow_291_fu_35690_p2 = (xor_ln895_453_fu_35684_p2 & p_Result_744_fu_35676_p3);

assign overflow_292_fu_35792_p2 = (xor_ln895_454_fu_35786_p2 & p_Result_746_fu_35778_p3);

assign overflow_293_fu_35894_p2 = (xor_ln895_455_fu_35888_p2 & p_Result_748_fu_35880_p3);

assign overflow_294_fu_35996_p2 = (xor_ln895_456_fu_35990_p2 & p_Result_750_fu_35982_p3);

assign overflow_295_fu_36098_p2 = (xor_ln895_457_fu_36092_p2 & p_Result_752_fu_36084_p3);

assign overflow_296_fu_36200_p2 = (xor_ln895_458_fu_36194_p2 & p_Result_754_fu_36186_p3);

assign overflow_297_fu_36302_p2 = (xor_ln895_459_fu_36296_p2 & p_Result_756_fu_36288_p3);

assign overflow_298_fu_36404_p2 = (xor_ln895_460_fu_36398_p2 & p_Result_758_fu_36390_p3);

assign overflow_299_fu_36506_p2 = (xor_ln895_461_fu_36500_p2 & p_Result_760_fu_36492_p3);

assign overflow_300_fu_36608_p2 = (xor_ln895_462_fu_36602_p2 & p_Result_762_fu_36594_p3);

assign overflow_301_fu_36710_p2 = (xor_ln895_463_fu_36704_p2 & p_Result_764_fu_36696_p3);

assign overflow_302_fu_36812_p2 = (xor_ln895_464_fu_36806_p2 & p_Result_766_fu_36798_p3);

assign overflow_303_fu_36914_p2 = (xor_ln895_465_fu_36908_p2 & p_Result_768_fu_36900_p3);

assign overflow_304_fu_37016_p2 = (xor_ln895_466_fu_37010_p2 & p_Result_770_fu_37002_p3);

assign overflow_305_fu_39442_p2 = (xor_ln895_467_fu_39436_p2 & p_Result_772_fu_39428_p3);

assign overflow_306_fu_39542_p2 = (xor_ln895_468_fu_39536_p2 & p_Result_774_fu_39528_p3);

assign overflow_307_fu_39642_p2 = (xor_ln895_469_fu_39636_p2 & p_Result_776_fu_39628_p3);

assign overflow_308_fu_39742_p2 = (xor_ln895_470_fu_39736_p2 & p_Result_778_fu_39728_p3);

assign overflow_309_fu_39842_p2 = (xor_ln895_471_fu_39836_p2 & p_Result_780_fu_39828_p3);

assign overflow_310_fu_39942_p2 = (xor_ln895_472_fu_39936_p2 & p_Result_782_fu_39928_p3);

assign overflow_311_fu_40042_p2 = (xor_ln895_473_fu_40036_p2 & p_Result_784_fu_40028_p3);

assign overflow_312_fu_40142_p2 = (xor_ln895_474_fu_40136_p2 & p_Result_786_fu_40128_p3);

assign overflow_313_fu_40242_p2 = (xor_ln895_475_fu_40236_p2 & p_Result_788_fu_40228_p3);

assign overflow_314_fu_40344_p2 = (xor_ln895_476_fu_40338_p2 & p_Result_790_fu_40330_p3);

assign overflow_315_fu_40446_p2 = (xor_ln895_477_fu_40440_p2 & p_Result_792_fu_40432_p3);

assign overflow_316_fu_40548_p2 = (xor_ln895_478_fu_40542_p2 & p_Result_794_fu_40534_p3);

assign overflow_317_fu_40650_p2 = (xor_ln895_479_fu_40644_p2 & p_Result_796_fu_40636_p3);

assign overflow_318_fu_40752_p2 = (xor_ln895_480_fu_40746_p2 & p_Result_798_fu_40738_p3);

assign overflow_319_fu_40854_p2 = (xor_ln895_481_fu_40848_p2 & p_Result_800_fu_40840_p3);

assign overflow_320_fu_40956_p2 = (xor_ln895_482_fu_40950_p2 & p_Result_802_fu_40942_p3);

assign overflow_321_fu_41058_p2 = (xor_ln895_483_fu_41052_p2 & p_Result_804_fu_41044_p3);

assign overflow_322_fu_41160_p2 = (xor_ln895_484_fu_41154_p2 & p_Result_806_fu_41146_p3);

assign overflow_fu_19040_p2 = (xor_ln895_243_fu_19035_p2 & or_ln895_fu_19030_p2);

assign p_Result_431_fu_20107_p3 = p_Val2_430_fu_20097_p2[32'd21];

assign p_Result_434_fu_20256_p3 = p_Val2_433_fu_20246_p2[32'd18];

assign p_Result_437_fu_20405_p3 = p_Val2_436_fu_20395_p2[32'd16];

assign p_Result_440_fu_20554_p3 = p_Val2_439_fu_20544_p2[32'd20];

assign p_Result_443_fu_20703_p3 = p_Val2_442_fu_20693_p2[32'd18];

assign p_Result_444_fu_18127_p3 = r_V_91_fu_18121_p2[32'd39];

assign p_Result_445_fu_18149_p3 = r_V_91_fu_18121_p2[32'd39];

assign p_Result_446_fu_18175_p3 = p_Val2_445_fu_18169_p2[32'd16];

assign p_Result_449_fu_20869_p3 = p_Val2_448_fu_20859_p2[32'd18];

assign p_Result_452_fu_21018_p3 = p_Val2_451_fu_21008_p2[32'd19];

assign p_Result_455_fu_21167_p3 = p_Val2_454_fu_21157_p2[32'd15];

assign p_Result_458_fu_21312_p3 = p_Val2_457_fu_21306_p2[32'd31];

assign p_Result_461_fu_21457_p3 = p_Val2_460_fu_21451_p2[32'd20];

assign p_Result_464_fu_21586_p3 = p_Val2_463_fu_21580_p2[32'd17];

assign p_Result_467_fu_21711_p3 = p_Val2_466_fu_21706_p2[32'd31];

assign p_Result_470_fu_21856_p3 = p_Val2_469_fu_21850_p2[32'd28];

assign p_Result_473_fu_21985_p3 = p_Val2_472_fu_21979_p2[32'd21];

assign p_Result_476_fu_22114_p3 = p_Val2_475_fu_22108_p2[32'd19];

assign p_Result_479_fu_22243_p3 = p_Val2_478_fu_22237_p2[32'd17];

assign p_Result_482_fu_22372_p3 = p_Val2_481_fu_22366_p2[32'd23];

assign p_Result_501_fu_22918_p3 = r_V_110_fu_22912_p2[32'd38];

assign p_Result_502_fu_22940_p3 = r_V_110_fu_22912_p2[32'd38];

assign p_Result_503_fu_22957_p3 = p_Val2_502_fu_22951_p2[32'd15];

assign p_Result_512_fu_26570_p3 = p_Val2_511_fu_26564_p2[32'd31];

assign p_Result_515_fu_26719_p3 = p_Val2_514_fu_26709_p2[32'd18];

assign p_Result_518_fu_26868_p3 = p_Val2_517_fu_26858_p2[32'd21];

assign p_Result_521_fu_27017_p3 = p_Val2_520_fu_27007_p2[32'd21];

assign p_Result_524_fu_27166_p3 = p_Val2_523_fu_27156_p2[32'd23];

assign p_Result_527_fu_27315_p3 = p_Val2_526_fu_27305_p2[32'd19];

assign p_Result_530_fu_27464_p3 = p_Val2_529_fu_27454_p2[32'd21];

assign p_Result_533_fu_27613_p3 = p_Val2_532_fu_27603_p2[32'd20];

assign p_Result_536_fu_27762_p3 = p_Val2_535_fu_27752_p2[32'd20];

assign p_Result_537_fu_27946_p3 = r_V_122_fu_27940_p2[32'd40];

assign p_Result_538_fu_27968_p3 = r_V_122_fu_27940_p2[32'd40];

assign p_Result_539_fu_27985_p3 = p_Val2_538_fu_27979_p2[32'd17];

assign p_Result_566_fu_32355_p3 = p_Val2_565_fu_32345_p2[32'd20];

assign p_Result_569_fu_32504_p3 = p_Val2_568_fu_32494_p2[32'd19];

assign p_Result_572_fu_32653_p3 = p_Val2_571_fu_32643_p2[32'd19];

assign p_Result_575_fu_32802_p3 = p_Val2_574_fu_32792_p2[32'd20];

assign p_Result_578_fu_32951_p3 = p_Val2_577_fu_32941_p2[32'd19];

assign p_Result_581_fu_33100_p3 = p_Val2_580_fu_33090_p2[32'd19];

assign p_Result_584_fu_33249_p3 = p_Val2_583_fu_33239_p2[32'd17];

assign p_Result_587_fu_33398_p3 = p_Val2_586_fu_33388_p2[32'd18];

assign p_Result_588_fu_29013_p3 = r_V_139_fu_29007_p2[32'd40];

assign p_Result_589_fu_29035_p3 = r_V_139_fu_29007_p2[32'd40];

assign p_Result_590_fu_29052_p3 = p_Val2_589_fu_29046_p2[32'd17];

assign p_Result_620_fu_38209_p3 = p_Val2_619_fu_38203_p2[32'd31];

assign p_Result_623_fu_38358_p3 = p_Val2_622_fu_38348_p2[32'd18];

assign p_Result_626_fu_38507_p3 = p_Val2_625_fu_38497_p2[32'd20];

assign p_Result_629_fu_38656_p3 = p_Val2_628_fu_38646_p2[32'd26];

assign p_Result_632_fu_38805_p3 = p_Val2_631_fu_38795_p2[32'd26];

assign p_Result_635_fu_38954_p3 = p_Val2_634_fu_38944_p2[32'd18];

assign p_Result_638_fu_39103_p3 = p_Val2_637_fu_39093_p2[32'd20];

assign p_Result_639_fu_34496_p3 = r_V_156_fu_34490_p2[32'd35];

assign p_Result_640_fu_34518_p3 = r_V_156_fu_34490_p2[32'd35];

assign p_Result_641_fu_34544_p3 = p_Val2_640_fu_34538_p2[32'd12];

assign p_Result_644_fu_39269_p3 = p_Val2_643_fu_39259_p2[32'd26];

assign p_Result_645_fu_23632_p3 = ret_V_fu_23626_p2[32'd32];

assign p_Result_646_fu_23646_p3 = p_Val2_645_fu_23640_p2[32'd31];

assign p_Result_647_fu_23730_p3 = ret_V_81_fu_23724_p2[32'd32];

assign p_Result_648_fu_23744_p3 = p_Val2_647_fu_23738_p2[32'd31];

assign p_Result_649_fu_23828_p3 = ret_V_82_fu_23822_p2[32'd32];

assign p_Result_650_fu_23842_p3 = p_Val2_649_fu_23836_p2[32'd31];

assign p_Result_651_fu_23926_p3 = ret_V_83_fu_23920_p2[32'd32];

assign p_Result_652_fu_23940_p3 = p_Val2_651_fu_23934_p2[32'd31];

assign p_Result_653_fu_24024_p3 = ret_V_84_fu_24018_p2[32'd32];

assign p_Result_654_fu_24038_p3 = p_Val2_653_fu_24032_p2[32'd31];

assign p_Result_655_fu_24122_p3 = ret_V_85_fu_24116_p2[32'd32];

assign p_Result_656_fu_24136_p3 = p_Val2_655_fu_24130_p2[32'd31];

assign p_Result_657_fu_24220_p3 = ret_V_86_fu_24214_p2[32'd32];

assign p_Result_658_fu_24234_p3 = p_Val2_657_fu_24228_p2[32'd31];

assign p_Result_659_fu_24318_p3 = ret_V_87_fu_24312_p2[32'd32];

assign p_Result_660_fu_24332_p3 = p_Val2_659_fu_24326_p2[32'd31];

assign p_Result_661_fu_24416_p3 = ret_V_88_fu_24410_p2[32'd32];

assign p_Result_662_fu_24430_p3 = p_Val2_661_fu_24424_p2[32'd31];

assign p_Result_663_fu_24518_p3 = ret_V_89_fu_24512_p2[32'd32];

assign p_Result_664_fu_24532_p3 = p_Val2_663_fu_24526_p2[32'd31];

assign p_Result_665_fu_24620_p3 = ret_V_90_fu_24614_p2[32'd32];

assign p_Result_666_fu_24634_p3 = p_Val2_665_fu_24628_p2[32'd31];

assign p_Result_667_fu_24722_p3 = ret_V_91_fu_24716_p2[32'd32];

assign p_Result_668_fu_24736_p3 = p_Val2_667_fu_24730_p2[32'd31];

assign p_Result_669_fu_24824_p3 = ret_V_92_fu_24818_p2[32'd32];

assign p_Result_670_fu_24838_p3 = p_Val2_669_fu_24832_p2[32'd31];

assign p_Result_671_fu_24926_p3 = ret_V_93_fu_24920_p2[32'd32];

assign p_Result_672_fu_24940_p3 = p_Val2_671_fu_24934_p2[32'd31];

assign p_Result_673_fu_25028_p3 = ret_V_94_fu_25022_p2[32'd32];

assign p_Result_674_fu_25042_p3 = p_Val2_673_fu_25036_p2[32'd31];

assign p_Result_675_fu_25130_p3 = ret_V_95_fu_25124_p2[32'd32];

assign p_Result_676_fu_25144_p3 = p_Val2_675_fu_25138_p2[32'd31];

assign p_Result_677_fu_25232_p3 = ret_V_96_fu_25226_p2[32'd32];

assign p_Result_678_fu_25246_p3 = p_Val2_677_fu_25240_p2[32'd31];

assign p_Result_679_fu_25334_p3 = ret_V_97_fu_25328_p2[32'd32];

assign p_Result_680_fu_25348_p3 = p_Val2_679_fu_25342_p2[32'd31];

assign p_Result_681_fu_29196_p3 = ret_V_98_fu_29190_p2[32'd32];

assign p_Result_682_fu_29208_p3 = p_Val2_681_fu_29204_p2[32'd31];

assign p_Result_683_fu_29295_p3 = ret_V_99_fu_29289_p2[32'd32];

assign p_Result_684_fu_29308_p3 = p_Val2_683_fu_29303_p2[32'd31];

assign p_Result_685_fu_29395_p3 = ret_V_100_fu_29389_p2[32'd32];

assign p_Result_686_fu_29408_p3 = p_Val2_685_fu_29403_p2[32'd31];

assign p_Result_687_fu_29494_p3 = ret_V_101_fu_29488_p2[32'd32];

assign p_Result_688_fu_29506_p3 = p_Val2_687_fu_29502_p2[32'd31];

assign p_Result_689_fu_29593_p3 = ret_V_102_fu_29587_p2[32'd32];

assign p_Result_690_fu_29606_p3 = p_Val2_689_fu_29601_p2[32'd31];

assign p_Result_691_fu_29693_p3 = ret_V_103_fu_29687_p2[32'd32];

assign p_Result_692_fu_29706_p3 = p_Val2_691_fu_29701_p2[32'd31];

assign p_Result_693_fu_29793_p3 = ret_V_104_fu_29787_p2[32'd32];

assign p_Result_694_fu_29806_p3 = p_Val2_693_fu_29801_p2[32'd31];

assign p_Result_695_fu_29893_p3 = ret_V_105_fu_29887_p2[32'd32];

assign p_Result_696_fu_29906_p3 = p_Val2_695_fu_29901_p2[32'd31];

assign p_Result_697_fu_29993_p3 = ret_V_106_fu_29987_p2[32'd32];

assign p_Result_698_fu_30006_p3 = p_Val2_697_fu_30001_p2[32'd31];

assign p_Result_699_fu_30094_p3 = ret_V_107_fu_30088_p2[32'd32];

assign p_Result_700_fu_30108_p3 = p_Val2_699_fu_30102_p2[32'd31];

assign p_Result_701_fu_30196_p3 = ret_V_108_fu_30190_p2[32'd32];

assign p_Result_702_fu_30210_p3 = p_Val2_701_fu_30204_p2[32'd31];

assign p_Result_703_fu_30298_p3 = ret_V_109_fu_30292_p2[32'd32];

assign p_Result_704_fu_30312_p3 = p_Val2_703_fu_30306_p2[32'd31];

assign p_Result_705_fu_30400_p3 = ret_V_110_fu_30394_p2[32'd32];

assign p_Result_706_fu_30414_p3 = p_Val2_705_fu_30408_p2[32'd31];

assign p_Result_707_fu_30502_p3 = ret_V_111_fu_30496_p2[32'd32];

assign p_Result_708_fu_30516_p3 = p_Val2_707_fu_30510_p2[32'd31];

assign p_Result_709_fu_30604_p3 = ret_V_112_fu_30598_p2[32'd32];

assign p_Result_710_fu_30618_p3 = p_Val2_709_fu_30612_p2[32'd31];

assign p_Result_711_fu_30706_p3 = ret_V_113_fu_30700_p2[32'd32];

assign p_Result_712_fu_30720_p3 = p_Val2_711_fu_30714_p2[32'd31];

assign p_Result_713_fu_30808_p3 = ret_V_114_fu_30802_p2[32'd32];

assign p_Result_714_fu_30822_p3 = p_Val2_713_fu_30816_p2[32'd31];

assign p_Result_715_fu_30910_p3 = ret_V_115_fu_30904_p2[32'd32];

assign p_Result_716_fu_30924_p3 = p_Val2_715_fu_30918_p2[32'd31];

assign p_Result_735_fu_35254_p3 = ret_V_125_fu_35248_p2[32'd32];

assign p_Result_736_fu_35268_p3 = p_Val2_735_fu_35262_p2[32'd31];

assign p_Result_737_fu_35356_p3 = ret_V_126_fu_35350_p2[32'd32];

assign p_Result_738_fu_35370_p3 = p_Val2_737_fu_35364_p2[32'd31];

assign p_Result_739_fu_35458_p3 = ret_V_127_fu_35452_p2[32'd32];

assign p_Result_740_fu_35472_p3 = p_Val2_739_fu_35466_p2[32'd31];

assign p_Result_741_fu_35560_p3 = ret_V_128_fu_35554_p2[32'd32];

assign p_Result_742_fu_35574_p3 = p_Val2_741_fu_35568_p2[32'd31];

assign p_Result_743_fu_35662_p3 = ret_V_129_fu_35656_p2[32'd32];

assign p_Result_744_fu_35676_p3 = p_Val2_743_fu_35670_p2[32'd31];

assign p_Result_745_fu_35764_p3 = ret_V_130_fu_35758_p2[32'd32];

assign p_Result_746_fu_35778_p3 = p_Val2_745_fu_35772_p2[32'd31];

assign p_Result_747_fu_35866_p3 = ret_V_131_fu_35860_p2[32'd32];

assign p_Result_748_fu_35880_p3 = p_Val2_747_fu_35874_p2[32'd31];

assign p_Result_749_fu_35968_p3 = ret_V_132_fu_35962_p2[32'd32];

assign p_Result_750_fu_35982_p3 = p_Val2_749_fu_35976_p2[32'd31];

assign p_Result_751_fu_36070_p3 = ret_V_133_fu_36064_p2[32'd32];

assign p_Result_752_fu_36084_p3 = p_Val2_751_fu_36078_p2[32'd31];

assign p_Result_753_fu_36172_p3 = ret_V_134_fu_36166_p2[32'd32];

assign p_Result_754_fu_36186_p3 = p_Val2_753_fu_36180_p2[32'd31];

assign p_Result_755_fu_36274_p3 = ret_V_135_fu_36268_p2[32'd32];

assign p_Result_756_fu_36288_p3 = p_Val2_755_fu_36282_p2[32'd31];

assign p_Result_757_fu_36376_p3 = ret_V_136_fu_36370_p2[32'd32];

assign p_Result_758_fu_36390_p3 = p_Val2_757_fu_36384_p2[32'd31];

assign p_Result_759_fu_36478_p3 = ret_V_137_fu_36472_p2[32'd32];

assign p_Result_760_fu_36492_p3 = p_Val2_759_fu_36486_p2[32'd31];

assign p_Result_761_fu_36580_p3 = ret_V_138_fu_36574_p2[32'd32];

assign p_Result_762_fu_36594_p3 = p_Val2_761_fu_36588_p2[32'd31];

assign p_Result_763_fu_36682_p3 = ret_V_139_fu_36676_p2[32'd32];

assign p_Result_764_fu_36696_p3 = p_Val2_763_fu_36690_p2[32'd31];

assign p_Result_765_fu_36784_p3 = ret_V_140_fu_36778_p2[32'd32];

assign p_Result_766_fu_36798_p3 = p_Val2_765_fu_36792_p2[32'd31];

assign p_Result_767_fu_36886_p3 = ret_V_141_fu_36880_p2[32'd32];

assign p_Result_768_fu_36900_p3 = p_Val2_767_fu_36894_p2[32'd31];

assign p_Result_769_fu_36988_p3 = ret_V_142_fu_36982_p2[32'd32];

assign p_Result_770_fu_37002_p3 = p_Val2_769_fu_36996_p2[32'd31];

assign p_Result_771_fu_39415_p3 = ret_V_143_fu_39409_p2[32'd32];

assign p_Result_772_fu_39428_p3 = p_Val2_771_fu_39423_p2[32'd31];

assign p_Result_773_fu_39515_p3 = ret_V_144_fu_39509_p2[32'd32];

assign p_Result_774_fu_39528_p3 = p_Val2_773_fu_39523_p2[32'd31];

assign p_Result_775_fu_39615_p3 = ret_V_145_fu_39609_p2[32'd32];

assign p_Result_776_fu_39628_p3 = p_Val2_775_fu_39623_p2[32'd31];

assign p_Result_777_fu_39715_p3 = ret_V_146_fu_39709_p2[32'd32];

assign p_Result_778_fu_39728_p3 = p_Val2_777_fu_39723_p2[32'd31];

assign p_Result_779_fu_39815_p3 = ret_V_147_fu_39809_p2[32'd32];

assign p_Result_780_fu_39828_p3 = p_Val2_779_fu_39823_p2[32'd31];

assign p_Result_781_fu_39915_p3 = ret_V_148_fu_39909_p2[32'd32];

assign p_Result_782_fu_39928_p3 = p_Val2_781_fu_39923_p2[32'd31];

assign p_Result_783_fu_40015_p3 = ret_V_149_fu_40009_p2[32'd32];

assign p_Result_784_fu_40028_p3 = p_Val2_783_fu_40023_p2[32'd31];

assign p_Result_785_fu_40115_p3 = ret_V_150_fu_40109_p2[32'd32];

assign p_Result_786_fu_40128_p3 = p_Val2_785_fu_40123_p2[32'd31];

assign p_Result_787_fu_40215_p3 = ret_V_151_fu_40209_p2[32'd32];

assign p_Result_788_fu_40228_p3 = p_Val2_787_fu_40223_p2[32'd31];

assign p_Result_789_fu_40316_p3 = ret_V_152_fu_40310_p2[32'd32];

assign p_Result_790_fu_40330_p3 = p_Val2_789_fu_40324_p2[32'd31];

assign p_Result_791_fu_40418_p3 = ret_V_153_fu_40412_p2[32'd32];

assign p_Result_792_fu_40432_p3 = p_Val2_791_fu_40426_p2[32'd31];

assign p_Result_793_fu_40520_p3 = ret_V_154_fu_40514_p2[32'd32];

assign p_Result_794_fu_40534_p3 = p_Val2_793_fu_40528_p2[32'd31];

assign p_Result_795_fu_40622_p3 = ret_V_155_fu_40616_p2[32'd32];

assign p_Result_796_fu_40636_p3 = p_Val2_795_fu_40630_p2[32'd31];

assign p_Result_797_fu_40724_p3 = ret_V_156_fu_40718_p2[32'd32];

assign p_Result_798_fu_40738_p3 = p_Val2_797_fu_40732_p2[32'd31];

assign p_Result_799_fu_40826_p3 = ret_V_157_fu_40820_p2[32'd32];

assign p_Result_800_fu_40840_p3 = p_Val2_799_fu_40834_p2[32'd31];

assign p_Result_801_fu_40928_p3 = ret_V_158_fu_40922_p2[32'd32];

assign p_Result_802_fu_40942_p3 = p_Val2_801_fu_40936_p2[32'd31];

assign p_Result_803_fu_41030_p3 = ret_V_159_fu_41024_p2[32'd32];

assign p_Result_804_fu_41044_p3 = p_Val2_803_fu_41038_p2[32'd31];

assign p_Result_805_fu_41132_p3 = ret_V_160_fu_41126_p2[32'd32];

assign p_Result_806_fu_41146_p3 = p_Val2_805_fu_41140_p2[32'd31];

assign p_Val2_402_fu_17281_p4 = {{r_V_fu_536_p2[41:24]}};

assign p_Val2_403_fu_17315_p2 = ($signed(zext_ln377_fu_17311_p1) + $signed(sext_ln823_fu_17291_p1));

assign p_Val2_405_fu_17345_p4 = {{r_V_78_fu_527_p2[42:24]}};

assign p_Val2_406_fu_17379_p2 = ($signed(zext_ln377_81_fu_17375_p1) + $signed(sext_ln823_78_fu_17355_p1));

assign p_Val2_408_fu_17409_p4 = {{r_V_79_fu_484_p2[43:24]}};

assign p_Val2_409_fu_17443_p2 = ($signed(zext_ln377_82_fu_17439_p1) + $signed(sext_ln823_79_fu_17419_p1));

assign p_Val2_411_fu_17473_p4 = {{r_V_80_fu_509_p2[41:24]}};

assign p_Val2_412_fu_17507_p2 = ($signed(zext_ln377_83_fu_17503_p1) + $signed(sext_ln823_80_fu_17483_p1));

assign p_Val2_414_fu_17537_p4 = {{r_V_81_fu_489_p2[41:24]}};

assign p_Val2_415_fu_17571_p2 = ($signed(zext_ln377_84_fu_17567_p1) + $signed(sext_ln823_81_fu_17547_p1));

assign p_Val2_417_fu_17601_p4 = {{r_V_82_fu_497_p2[43:24]}};

assign p_Val2_418_fu_17635_p2 = ($signed(zext_ln377_85_fu_17631_p1) + $signed(sext_ln823_82_fu_17611_p1));

assign p_Val2_420_fu_17665_p4 = {{r_V_83_fu_507_p2[44:24]}};

assign p_Val2_421_fu_17699_p2 = ($signed(zext_ln377_86_fu_17695_p1) + $signed(sext_ln823_83_fu_17675_p1));

assign p_Val2_423_fu_17729_p4 = {{r_V_84_fu_494_p2[39:24]}};

assign p_Val2_424_fu_17763_p2 = ($signed(zext_ln377_87_fu_17759_p1) + $signed(sext_ln823_84_fu_17739_p1));

assign p_Val2_426_fu_17793_p4 = {{r_V_85_fu_495_p2[42:24]}};

assign p_Val2_427_fu_17827_p2 = ($signed(zext_ln377_88_fu_17823_p1) + $signed(sext_ln823_85_fu_17803_p1));

assign p_Val2_430_fu_20097_p2 = ($signed(zext_ln377_89_fu_20094_p1) + $signed(sext_ln823_86_fu_20091_p1));

assign p_Val2_433_fu_20246_p2 = ($signed(zext_ln377_90_fu_20243_p1) + $signed(sext_ln823_87_fu_20240_p1));

assign p_Val2_436_fu_20395_p2 = ($signed(zext_ln377_91_fu_20392_p1) + $signed(sext_ln823_88_fu_20389_p1));

assign p_Val2_439_fu_20544_p2 = ($signed(zext_ln377_92_fu_20541_p1) + $signed(sext_ln823_89_fu_20538_p1));

assign p_Val2_442_fu_20693_p2 = ($signed(zext_ln377_93_fu_20690_p1) + $signed(sext_ln823_90_fu_20687_p1));

assign p_Val2_444_fu_18135_p4 = {{r_V_91_fu_18121_p2[39:24]}};

assign p_Val2_445_fu_18169_p2 = ($signed(zext_ln377_94_fu_18165_p1) + $signed(sext_ln823_91_fu_18145_p1));

assign p_Val2_448_fu_20859_p2 = ($signed(zext_ln377_95_fu_20856_p1) + $signed(sext_ln823_92_fu_20853_p1));

assign p_Val2_451_fu_21008_p2 = ($signed(zext_ln377_96_fu_21005_p1) + $signed(sext_ln823_93_fu_21002_p1));

assign p_Val2_454_fu_21157_p2 = ($signed(zext_ln377_97_fu_21154_p1) + $signed(sext_ln823_94_fu_21151_p1));

assign p_Val2_457_fu_21306_p2 = ($signed(zext_ln377_98_fu_21303_p1) + $signed(sext_ln818_fu_21300_p1));

assign p_Val2_460_fu_21451_p2 = ($signed(zext_ln377_99_fu_21448_p1) + $signed(sext_ln823_95_fu_21445_p1));

assign p_Val2_463_fu_21580_p2 = ($signed(zext_ln377_100_fu_21577_p1) + $signed(sext_ln823_96_fu_21574_p1));

assign p_Val2_466_fu_21706_p2 = (zext_ln377_101_fu_21703_p1 + p_Val2_465_reg_41952);

assign p_Val2_469_fu_21850_p2 = ($signed(zext_ln377_102_fu_21847_p1) + $signed(sext_ln823_97_fu_21844_p1));

assign p_Val2_472_fu_21979_p2 = ($signed(zext_ln377_103_fu_21976_p1) + $signed(sext_ln823_98_fu_21973_p1));

assign p_Val2_475_fu_22108_p2 = ($signed(zext_ln377_104_fu_22105_p1) + $signed(sext_ln823_99_fu_22102_p1));

assign p_Val2_478_fu_22237_p2 = ($signed(zext_ln377_105_fu_22234_p1) + $signed(sext_ln823_100_fu_22231_p1));

assign p_Val2_481_fu_22366_p2 = ($signed(zext_ln377_106_fu_22363_p1) + $signed(sext_ln823_101_fu_22360_p1));

assign p_Val2_483_fu_22514_p4 = {{r_V_104_fu_466_p2[41:24]}};

assign p_Val2_484_fu_22548_p2 = ($signed(zext_ln377_107_fu_22544_p1) + $signed(sext_ln823_102_fu_22524_p1));

assign p_Val2_486_fu_22578_p4 = {{r_V_105_fu_539_p2[42:24]}};

assign p_Val2_487_fu_22612_p2 = ($signed(zext_ln377_108_fu_22608_p1) + $signed(sext_ln823_103_fu_22588_p1));

assign p_Val2_489_fu_22642_p4 = {{r_V_106_fu_512_p2[41:24]}};

assign p_Val2_490_fu_22676_p2 = ($signed(zext_ln377_109_fu_22672_p1) + $signed(sext_ln823_104_fu_22652_p1));

assign p_Val2_492_fu_22706_p4 = {{r_V_107_fu_463_p2[42:24]}};

assign p_Val2_493_fu_22740_p2 = ($signed(zext_ln377_110_fu_22736_p1) + $signed(sext_ln823_105_fu_22716_p1));

assign p_Val2_495_fu_22770_p4 = {{r_V_108_fu_529_p2[43:24]}};

assign p_Val2_496_fu_22804_p2 = ($signed(zext_ln377_111_fu_22800_p1) + $signed(sext_ln823_106_fu_22780_p1));

assign p_Val2_498_fu_22834_p4 = {{r_V_109_fu_485_p2[41:24]}};

assign p_Val2_499_fu_22868_p2 = ($signed(zext_ln377_112_fu_22864_p1) + $signed(sext_ln823_107_fu_22844_p1));

assign p_Val2_501_fu_22926_p4 = {{r_V_110_fu_22912_p2[38:24]}};

assign p_Val2_502_fu_22951_p2 = ($signed(zext_ln377_113_fu_22948_p1) + $signed(sext_ln823_108_fu_22936_p1));

assign p_Val2_504_fu_23097_p4 = {{r_V_111_fu_526_p2[43:24]}};

assign p_Val2_505_fu_23131_p2 = ($signed(zext_ln377_114_fu_23127_p1) + $signed(sext_ln823_109_fu_23107_p1));

assign p_Val2_507_fu_23161_p4 = {{r_V_112_fu_471_p2[42:24]}};

assign p_Val2_508_fu_23195_p2 = ($signed(zext_ln377_115_fu_23191_p1) + $signed(sext_ln823_110_fu_23171_p1));

assign p_Val2_511_fu_26564_p2 = ($signed(zext_ln377_116_fu_26561_p1) + $signed(sext_ln818_1_fu_26558_p1));

assign p_Val2_514_fu_26709_p2 = ($signed(zext_ln377_117_fu_26706_p1) + $signed(sext_ln823_111_fu_26703_p1));

assign p_Val2_517_fu_26858_p2 = ($signed(zext_ln377_118_fu_26855_p1) + $signed(sext_ln823_112_fu_26852_p1));

assign p_Val2_520_fu_27007_p2 = ($signed(zext_ln377_119_fu_27004_p1) + $signed(sext_ln823_113_fu_27001_p1));

assign p_Val2_523_fu_27156_p2 = ($signed(zext_ln377_120_fu_27153_p1) + $signed(sext_ln823_114_fu_27150_p1));

assign p_Val2_526_fu_27305_p2 = ($signed(zext_ln377_121_fu_27302_p1) + $signed(sext_ln823_115_fu_27299_p1));

assign p_Val2_529_fu_27454_p2 = ($signed(zext_ln377_122_fu_27451_p1) + $signed(sext_ln823_116_fu_27448_p1));

assign p_Val2_532_fu_27603_p2 = ($signed(zext_ln377_123_fu_27600_p1) + $signed(sext_ln823_117_fu_27597_p1));

assign p_Val2_535_fu_27752_p2 = ($signed(zext_ln377_124_fu_27749_p1) + $signed(sext_ln823_118_fu_27746_p1));

assign p_Val2_537_fu_27954_p4 = {{r_V_122_fu_27940_p2[40:24]}};

assign p_Val2_538_fu_27979_p2 = ($signed(zext_ln377_125_fu_27976_p1) + $signed(sext_ln823_119_fu_27964_p1));

assign p_Val2_540_fu_28125_p4 = {{r_V_123_fu_472_p2[42:24]}};

assign p_Val2_541_fu_28159_p2 = ($signed(zext_ln377_126_fu_28155_p1) + $signed(sext_ln823_120_fu_28135_p1));

assign p_Val2_543_fu_28189_p4 = {{r_V_124_fu_462_p2[43:24]}};

assign p_Val2_544_fu_28223_p2 = ($signed(zext_ln377_127_fu_28219_p1) + $signed(sext_ln823_121_fu_28199_p1));

assign p_Val2_546_fu_28253_p4 = {{r_V_125_fu_510_p2[42:24]}};

assign p_Val2_547_fu_28287_p2 = ($signed(zext_ln377_128_fu_28283_p1) + $signed(sext_ln823_122_fu_28263_p1));

assign p_Val2_549_fu_28317_p4 = {{r_V_126_fu_515_p2[43:24]}};

assign p_Val2_550_fu_28351_p2 = ($signed(zext_ln377_129_fu_28347_p1) + $signed(sext_ln823_123_fu_28327_p1));

assign p_Val2_552_fu_28381_p4 = {{r_V_127_fu_479_p2[42:24]}};

assign p_Val2_553_fu_28415_p2 = ($signed(zext_ln377_130_fu_28411_p1) + $signed(sext_ln823_124_fu_28391_p1));

assign p_Val2_555_fu_28445_p4 = {{r_V_128_fu_513_p2[44:24]}};

assign p_Val2_556_fu_28479_p2 = ($signed(zext_ln377_131_fu_28475_p1) + $signed(sext_ln823_125_fu_28455_p1));

assign p_Val2_558_fu_28509_p4 = {{r_V_129_fu_521_p2[39:24]}};

assign p_Val2_559_fu_28543_p2 = ($signed(zext_ln377_132_fu_28539_p1) + $signed(sext_ln823_126_fu_28519_p1));

assign p_Val2_561_fu_28573_p4 = {{r_V_130_fu_491_p2[41:24]}};

assign p_Val2_562_fu_28607_p2 = ($signed(zext_ln377_133_fu_28603_p1) + $signed(sext_ln823_127_fu_28583_p1));

assign p_Val2_565_fu_32345_p2 = ($signed(zext_ln377_134_fu_32342_p1) + $signed(sext_ln823_128_fu_32339_p1));

assign p_Val2_568_fu_32494_p2 = ($signed(zext_ln377_135_fu_32491_p1) + $signed(sext_ln823_129_fu_32488_p1));

assign p_Val2_571_fu_32643_p2 = ($signed(zext_ln377_136_fu_32640_p1) + $signed(sext_ln823_130_fu_32637_p1));

assign p_Val2_574_fu_32792_p2 = ($signed(zext_ln377_137_fu_32789_p1) + $signed(sext_ln823_131_fu_32786_p1));

assign p_Val2_577_fu_32941_p2 = ($signed(zext_ln377_138_fu_32938_p1) + $signed(sext_ln823_132_fu_32935_p1));

assign p_Val2_580_fu_33090_p2 = ($signed(zext_ln377_139_fu_33087_p1) + $signed(sext_ln823_133_fu_33084_p1));

assign p_Val2_583_fu_33239_p2 = ($signed(zext_ln377_140_fu_33236_p1) + $signed(sext_ln823_134_fu_33233_p1));

assign p_Val2_586_fu_33388_p2 = ($signed(zext_ln377_141_fu_33385_p1) + $signed(sext_ln823_135_fu_33382_p1));

assign p_Val2_588_fu_29021_p4 = {{r_V_139_fu_29007_p2[40:24]}};

assign p_Val2_589_fu_29046_p2 = ($signed(zext_ln377_142_fu_29043_p1) + $signed(sext_ln823_136_fu_29031_p1));

assign p_Val2_591_fu_33580_p4 = {{r_V_140_fu_481_p2[54:24]}};

assign p_Val2_592_fu_33614_p2 = ($signed(zext_ln377_143_fu_33610_p1) + $signed(sext_ln818_2_fu_33590_p1));

assign p_Val2_594_fu_33644_p4 = {{r_V_141_fu_541_p2[43:24]}};

assign p_Val2_595_fu_33678_p2 = ($signed(zext_ln377_144_fu_33674_p1) + $signed(sext_ln823_137_fu_33654_p1));

assign p_Val2_597_fu_33708_p4 = {{r_V_142_fu_492_p2[42:24]}};

assign p_Val2_598_fu_33742_p2 = ($signed(zext_ln377_145_fu_33738_p1) + $signed(sext_ln823_138_fu_33718_p1));

assign p_Val2_600_fu_33772_p4 = {{r_V_143_fu_540_p2[49:24]}};

assign p_Val2_601_fu_33806_p2 = ($signed(zext_ln377_146_fu_33802_p1) + $signed(sext_ln823_139_fu_33782_p1));

assign p_Val2_603_fu_33836_p4 = {{r_V_144_fu_490_p2[48:24]}};

assign p_Val2_604_fu_33870_p2 = ($signed(zext_ln377_147_fu_33866_p1) + $signed(sext_ln823_140_fu_33846_p1));

assign p_Val2_606_fu_33900_p4 = {{r_V_145_fu_476_p2[43:24]}};

assign p_Val2_607_fu_33934_p2 = ($signed(zext_ln377_148_fu_33930_p1) + $signed(sext_ln823_141_fu_33910_p1));

assign p_Val2_609_fu_33964_p4 = {{r_V_146_fu_514_p2[43:24]}};

assign p_Val2_610_fu_33998_p2 = ($signed(zext_ln377_149_fu_33994_p1) + $signed(sext_ln823_142_fu_33974_p1));

assign p_Val2_612_fu_34028_p4 = {{r_V_147_fu_508_p2[43:24]}};

assign p_Val2_613_fu_34062_p2 = ($signed(zext_ln377_150_fu_34058_p1) + $signed(sext_ln823_143_fu_34038_p1));

assign p_Val2_615_fu_34092_p4 = {{r_V_148_fu_518_p2[48:24]}};

assign p_Val2_616_fu_34126_p2 = ($signed(zext_ln377_151_fu_34122_p1) + $signed(sext_ln823_144_fu_34102_p1));

assign p_Val2_619_fu_38203_p2 = ($signed(zext_ln377_152_fu_38200_p1) + $signed(sext_ln818_3_fu_38197_p1));

assign p_Val2_622_fu_38348_p2 = ($signed(zext_ln377_153_fu_38345_p1) + $signed(sext_ln823_145_fu_38342_p1));

assign p_Val2_625_fu_38497_p2 = ($signed(zext_ln377_154_fu_38494_p1) + $signed(sext_ln823_146_fu_38491_p1));

assign p_Val2_628_fu_38646_p2 = ($signed(zext_ln377_155_fu_38643_p1) + $signed(sext_ln823_147_fu_38640_p1));

assign p_Val2_631_fu_38795_p2 = ($signed(zext_ln377_156_fu_38792_p1) + $signed(sext_ln823_148_fu_38789_p1));

assign p_Val2_634_fu_38944_p2 = ($signed(zext_ln377_157_fu_38941_p1) + $signed(sext_ln823_149_fu_38938_p1));

assign p_Val2_637_fu_39093_p2 = ($signed(zext_ln377_158_fu_39090_p1) + $signed(sext_ln823_150_fu_39087_p1));

assign p_Val2_639_fu_34504_p4 = {{r_V_156_fu_34490_p2[35:24]}};

assign p_Val2_640_fu_34538_p2 = ($signed(zext_ln377_159_fu_34534_p1) + $signed(sext_ln823_151_fu_34514_p1));

assign p_Val2_643_fu_39259_p2 = ($signed(zext_ln377_160_fu_39256_p1) + $signed(sext_ln823_152_fu_39253_p1));

assign p_Val2_645_fu_23640_p2 = ($signed(rhs_fu_19083_p3) + $signed(32'd5264183));

assign p_Val2_647_fu_23738_p2 = ($signed(rhs_81_fu_19208_p3) + $signed(32'd4294918003));

assign p_Val2_649_fu_23836_p2 = ($signed(rhs_82_fu_19333_p3) + $signed(32'd4294373753));

assign p_Val2_651_fu_23934_p2 = ($signed(rhs_83_fu_19458_p3) + $signed(32'd4294962125));

assign p_Val2_653_fu_24032_p2 = ($signed(rhs_84_fu_19583_p3) + $signed(32'd6442053));

assign p_Val2_655_fu_24130_p2 = ($signed(rhs_85_fu_19708_p3) + $signed(32'd4294963189));

assign p_Val2_657_fu_24228_p2 = ($signed(rhs_86_fu_19833_p3) + $signed(32'd4294812477));

assign p_Val2_659_fu_24326_p2 = ($signed(rhs_87_fu_19958_p3) + $signed(32'd4294753504));

assign p_Val2_661_fu_24424_p2 = ($signed(rhs_88_fu_20083_p3) + $signed(32'd19328802));

assign p_Val2_663_fu_24526_p2 = ($signed(rhs_89_fu_20232_p3) + $signed(lhs_fu_23712_p3));

assign p_Val2_665_fu_24628_p2 = ($signed(rhs_90_fu_20381_p3) + $signed(lhs_72_fu_23810_p3));

assign p_Val2_667_fu_24730_p2 = ($signed(rhs_91_fu_20530_p3) + $signed(lhs_73_fu_23908_p3));

assign p_Val2_669_fu_24832_p2 = ($signed(rhs_92_fu_20679_p3) + $signed(lhs_74_fu_24006_p3));

assign p_Val2_671_fu_24934_p2 = ($signed(rhs_93_fu_20828_p3) + $signed(lhs_75_fu_24104_p3));

assign p_Val2_673_fu_25036_p2 = ($signed(rhs_94_fu_20846_p3) + $signed(lhs_76_fu_24202_p3));

assign p_Val2_675_fu_25138_p2 = ($signed(rhs_95_fu_20994_p3) + $signed(lhs_77_fu_24300_p3));

assign p_Val2_677_fu_25240_p2 = ($signed(rhs_96_fu_21143_p3) + $signed(lhs_78_fu_24398_p3));

assign p_Val2_679_fu_25342_p2 = ($signed(rhs_97_fu_21292_p3) + $signed(lhs_79_fu_24496_p3));

assign p_Val2_681_fu_29204_p2 = ($signed(rhs_98_reg_42135) + $signed(lhs_80_reg_42776));

assign p_Val2_683_fu_29303_p2 = ($signed(rhs_99_fu_25432_p3) + $signed(lhs_81_reg_42782));

assign p_Val2_685_fu_29403_p2 = ($signed(rhs_100_fu_25449_p3) + $signed(lhs_82_reg_42788));

assign p_Val2_687_fu_29502_p2 = ($signed(rhs_101_reg_42171) + $signed(lhs_83_reg_42794));

assign p_Val2_689_fu_29601_p2 = ($signed(rhs_102_fu_25466_p3) + $signed(lhs_84_reg_42800));

assign p_Val2_691_fu_29701_p2 = ($signed(rhs_103_fu_25483_p3) + $signed(lhs_85_reg_42806));

assign p_Val2_693_fu_29801_p2 = ($signed(rhs_104_fu_25500_p3) + $signed(lhs_86_reg_42812));

assign p_Val2_695_fu_29901_p2 = ($signed(rhs_105_fu_25517_p3) + $signed(lhs_87_reg_42818));

assign p_Val2_697_fu_30001_p2 = ($signed(rhs_106_fu_25534_p3) + $signed(lhs_88_reg_42824));

assign p_Val2_699_fu_30102_p2 = ($signed(rhs_107_fu_25658_p3) + $signed(lhs_89_fu_29274_p3));

assign p_Val2_701_fu_30204_p2 = ($signed(rhs_108_fu_25783_p3) + $signed(lhs_90_fu_29374_p3));

assign p_Val2_703_fu_30306_p2 = ($signed(rhs_109_fu_25908_p3) + $signed(lhs_91_fu_29474_p3));

assign p_Val2_705_fu_30408_p2 = ($signed(rhs_110_fu_26033_p3) + $signed(lhs_92_fu_29572_p3));

assign p_Val2_707_fu_30510_p2 = ($signed(rhs_111_fu_26158_p3) + $signed(lhs_93_fu_29672_p3));

assign p_Val2_709_fu_30612_p2 = ($signed(rhs_112_fu_26283_p3) + $signed(lhs_94_fu_29772_p3));

assign p_Val2_711_fu_30714_p2 = ($signed(rhs_113_fu_26301_p3) + $signed(lhs_95_fu_29872_p3));

assign p_Val2_713_fu_30816_p2 = ($signed(rhs_114_fu_26425_p3) + $signed(lhs_96_fu_29972_p3));

assign p_Val2_715_fu_30918_p2 = ($signed(rhs_115_fu_26550_p3) + $signed(lhs_97_fu_30072_p3));

assign p_Val2_717_fu_31020_p2 = ($signed(rhs_116_fu_26695_p3) + $signed(lhs_98_fu_30174_p3));

assign p_Val2_719_fu_31056_p2 = ($signed(rhs_117_fu_26844_p3) + $signed(lhs_99_fu_30276_p3));

assign p_Val2_721_fu_31092_p2 = ($signed(rhs_118_fu_26993_p3) + $signed(lhs_100_fu_30378_p3));

assign p_Val2_723_fu_31128_p2 = ($signed(rhs_119_fu_27142_p3) + $signed(lhs_101_fu_30480_p3));

assign p_Val2_725_fu_31164_p2 = ($signed(rhs_120_fu_27291_p3) + $signed(lhs_102_fu_30582_p3));

assign p_Val2_727_fu_31200_p2 = ($signed(rhs_121_fu_27440_p3) + $signed(lhs_103_fu_30684_p3));

assign p_Val2_729_fu_31236_p2 = ($signed(rhs_122_fu_27589_p3) + $signed(lhs_104_fu_30786_p3));

assign p_Val2_731_fu_31272_p2 = ($signed(rhs_123_fu_27738_p3) + $signed(lhs_105_fu_30888_p3));

assign p_Val2_733_fu_31308_p2 = ($signed(rhs_124_fu_27887_p3) + $signed(lhs_106_fu_30990_p3));

assign p_Val2_735_fu_35262_p2 = ($signed(rhs_125_fu_31332_p3) + $signed(lhs_107_fu_34768_p3));

assign p_Val2_737_fu_35364_p2 = ($signed(rhs_126_fu_31456_p3) + $signed(lhs_108_fu_34826_p3));

assign p_Val2_739_fu_35466_p2 = ($signed(rhs_127_fu_31581_p3) + $signed(lhs_109_fu_34884_p3));

assign p_Val2_741_fu_35568_p2 = ($signed(rhs_128_fu_31706_p3) + $signed(lhs_110_fu_34942_p3));

assign p_Val2_743_fu_35670_p2 = ($signed(rhs_129_fu_31831_p3) + $signed(lhs_111_fu_35000_p3));

assign p_Val2_745_fu_35772_p2 = ($signed(rhs_130_fu_31956_p3) + $signed(lhs_112_fu_35058_p3));

assign p_Val2_747_fu_35874_p2 = ($signed(rhs_131_fu_32081_p3) + $signed(lhs_113_fu_35116_p3));

assign p_Val2_749_fu_35976_p2 = ($signed(rhs_132_fu_32206_p3) + $signed(lhs_114_fu_35174_p3));

assign p_Val2_751_fu_36078_p2 = ($signed(rhs_133_fu_32331_p3) + $signed(lhs_115_fu_35232_p3));

assign p_Val2_753_fu_36180_p2 = ($signed(rhs_134_fu_32480_p3) + $signed(lhs_116_fu_35334_p3));

assign p_Val2_755_fu_36282_p2 = ($signed(rhs_135_fu_32629_p3) + $signed(lhs_117_fu_35436_p3));

assign p_Val2_757_fu_36384_p2 = ($signed(rhs_136_fu_32778_p3) + $signed(lhs_118_fu_35538_p3));

assign p_Val2_759_fu_36486_p2 = ($signed(rhs_137_fu_32927_p3) + $signed(lhs_119_fu_35640_p3));

assign p_Val2_761_fu_36588_p2 = ($signed(rhs_138_fu_33076_p3) + $signed(lhs_120_fu_35742_p3));

assign p_Val2_763_fu_36690_p2 = ($signed(rhs_139_fu_33225_p3) + $signed(lhs_121_fu_35844_p3));

assign p_Val2_765_fu_36792_p2 = ($signed(rhs_140_fu_33374_p3) + $signed(lhs_122_fu_35946_p3));

assign p_Val2_767_fu_36894_p2 = ($signed(rhs_141_fu_33523_p3) + $signed(lhs_123_fu_36048_p3));

assign p_Val2_769_fu_36996_p2 = ($signed(rhs_142_fu_33541_p3) + $signed(lhs_124_fu_36150_p3));

assign p_Val2_771_fu_39423_p2 = ($signed(rhs_143_fu_37190_p3) + $signed(lhs_125_reg_44046));

assign p_Val2_773_fu_39523_p2 = ($signed(rhs_144_fu_37314_p3) + $signed(lhs_126_reg_44052));

assign p_Val2_775_fu_39623_p2 = ($signed(rhs_145_fu_37439_p3) + $signed(lhs_127_reg_44058));

assign p_Val2_777_fu_39723_p2 = ($signed(rhs_146_fu_37564_p3) + $signed(lhs_128_reg_44064));

assign p_Val2_779_fu_39823_p2 = ($signed(rhs_147_fu_37689_p3) + $signed(lhs_129_reg_44070));

assign p_Val2_781_fu_39923_p2 = ($signed(rhs_148_fu_37814_p3) + $signed(lhs_130_reg_44076));

assign p_Val2_783_fu_40023_p2 = ($signed(rhs_149_fu_37939_p3) + $signed(lhs_131_reg_44082));

assign p_Val2_785_fu_40123_p2 = ($signed(rhs_150_fu_38064_p3) + $signed(lhs_132_reg_44088));

assign p_Val2_787_fu_40223_p2 = ($signed(rhs_151_fu_38189_p3) + $signed(lhs_133_reg_44094));

assign p_Val2_789_fu_40324_p2 = ($signed(rhs_152_fu_38334_p3) + $signed(lhs_134_fu_39494_p3));

assign p_Val2_791_fu_40426_p2 = ($signed(rhs_153_fu_38483_p3) + $signed(lhs_135_fu_39594_p3));

assign p_Val2_793_fu_40528_p2 = ($signed(rhs_154_fu_38632_p3) + $signed(lhs_136_fu_39694_p3));

assign p_Val2_795_fu_40630_p2 = ($signed(rhs_155_fu_38781_p3) + $signed(lhs_137_fu_39794_p3));

assign p_Val2_797_fu_40732_p2 = ($signed(rhs_156_fu_38930_p3) + $signed(lhs_138_fu_39894_p3));

assign p_Val2_799_fu_40834_p2 = ($signed(rhs_157_fu_39079_p3) + $signed(lhs_139_fu_39994_p3));

assign p_Val2_801_fu_40936_p2 = ($signed(rhs_158_fu_39228_p3) + $signed(lhs_140_fu_40094_p3));

assign p_Val2_803_fu_41038_p2 = ($signed(rhs_159_fu_39246_p3) + $signed(lhs_141_fu_40194_p3));

assign p_Val2_805_fu_41140_p2 = ($signed(rhs_160_fu_39394_p3) + $signed(lhs_142_fu_40294_p3));

assign r_V_100_fu_534_p1 = 45'd35184372086677;

assign r_V_101_fu_478_p1 = 43'd952;

assign r_V_102_fu_474_p0 = sext_ln70_60_fu_18458_p1;

assign r_V_102_fu_474_p1 = 41'd223;

assign r_V_103_fu_469_p1 = 47'd140737488341606;

assign r_V_104_fu_466_p0 = sext_ln70_65_fu_22500_p1;

assign r_V_104_fu_466_p1 = 42'd4398046510603;

assign r_V_105_fu_539_p0 = sext_ln70_64_fu_22494_p1;

assign r_V_105_fu_539_p1 = 43'd8796093021532;

assign r_V_106_fu_512_p0 = sext_ln70_65_fu_22500_p1;

assign r_V_106_fu_512_p1 = 42'd4398046510837;

assign r_V_107_fu_463_p0 = sext_ln70_64_fu_22494_p1;

assign r_V_107_fu_463_p1 = 43'd8796093021284;

assign r_V_108_fu_529_p0 = sext_ln70_63_fu_22489_p1;

assign r_V_108_fu_529_p1 = 44'd1275;

assign r_V_109_fu_485_p0 = sext_ln70_65_fu_22500_p1;

assign r_V_109_fu_485_p1 = 42'd446;

assign r_V_110_fu_22912_p2 = ($signed(sext_ln1273_15_fu_22908_p1) - $signed(sext_ln1273_14_fu_22897_p1));

assign r_V_111_fu_526_p0 = sext_ln70_63_fu_22489_p1;

assign r_V_111_fu_526_p1 = 44'd2026;

assign r_V_112_fu_471_p0 = sext_ln70_64_fu_22494_p1;

assign r_V_112_fu_471_p1 = 43'd894;

assign r_V_113_fu_535_p1 = 55'd5944544;

assign r_V_114_fu_475_p1 = 42'd4398046510628;

assign r_V_115_fu_468_p0 = sext_ln70_69_fu_23230_p1;

assign r_V_115_fu_468_p1 = 45'd35184372086675;

assign r_V_116_fu_537_p0 = sext_ln70_69_fu_23230_p1;

assign r_V_116_fu_537_p1 = 45'd35184372086038;

assign r_V_117_fu_519_p1 = 47'd140737488342760;

assign r_V_118_fu_470_p1 = 43'd8796093021313;

assign r_V_119_fu_542_p0 = sext_ln70_69_fu_23230_p1;

assign r_V_119_fu_542_p1 = 45'd2798;

assign r_V_120_fu_520_p0 = sext_ln70_66_fu_23217_p1;

assign r_V_120_fu_520_p1 = 44'd1303;

assign r_V_121_fu_477_p0 = sext_ln70_66_fu_23217_p1;

assign r_V_121_fu_477_p1 = 44'd17592186042845;

assign r_V_122_fu_27940_p2 = ($signed(sext_ln1273_17_fu_27936_p1) - $signed(sext_ln1273_16_fu_27925_p1));

assign r_V_123_fu_472_p0 = sext_ln70_75_fu_27908_p1;

assign r_V_123_fu_472_p1 = 43'd845;

assign r_V_124_fu_462_p0 = sext_ln70_74_fu_27903_p1;

assign r_V_124_fu_462_p1 = 44'd1062;

assign r_V_125_fu_510_p0 = sext_ln70_75_fu_27908_p1;

assign r_V_125_fu_510_p1 = 43'd910;

assign r_V_126_fu_515_p0 = sext_ln70_74_fu_27903_p1;

assign r_V_126_fu_515_p1 = 44'd17592186043118;

assign r_V_127_fu_479_p0 = sext_ln70_75_fu_27908_p1;

assign r_V_127_fu_479_p1 = 43'd739;

assign r_V_128_fu_513_p1 = 45'd2091;

assign r_V_129_fu_521_p1 = 40'd67;

assign r_V_130_fu_491_p1 = 42'd4398046510833;

assign r_V_131_fu_506_p0 = sext_ln70_80_fu_28644_p1;

assign r_V_131_fu_506_p1 = 44'd17592186042909;

assign r_V_132_fu_533_p0 = sext_ln70_79_fu_28637_p1;

assign r_V_132_fu_533_p1 = 43'd8796093021483;

assign r_V_133_fu_486_p0 = sext_ln70_79_fu_28637_p1;

assign r_V_133_fu_486_p1 = 43'd778;

assign r_V_134_fu_525_p0 = sext_ln70_80_fu_28644_p1;

assign r_V_134_fu_525_p1 = 44'd17592186043029;

assign r_V_135_fu_496_p0 = sext_ln70_79_fu_28637_p1;

assign r_V_135_fu_496_p1 = 43'd595;

assign r_V_136_fu_500_p0 = sext_ln70_79_fu_28637_p1;

assign r_V_136_fu_500_p1 = 43'd8796093021222;

assign r_V_137_fu_464_p1 = 41'd2199023255368;

assign r_V_138_fu_528_p1 = 42'd280;

assign r_V_139_fu_29007_p2 = ($signed(sext_ln1273_19_fu_29003_p1) - $signed(sext_ln1273_18_fu_28992_p1));

assign r_V_140_fu_481_p1 = 55'd36028797011804136;

assign r_V_141_fu_541_p0 = sext_ln70_84_fu_33561_p1;

assign r_V_141_fu_541_p1 = 44'd17592186043027;

assign r_V_142_fu_492_p1 = 43'd8796093021404;

assign r_V_143_fu_540_p1 = 50'd1125899906763676;

assign r_V_144_fu_490_p0 = sext_ln70_81_fu_33548_p1;

assign r_V_144_fu_490_p1 = 49'd41389;

assign r_V_145_fu_476_p0 = sext_ln70_84_fu_33561_p1;

assign r_V_145_fu_476_p1 = 44'd17592186043363;

assign r_V_146_fu_514_p0 = sext_ln70_84_fu_33561_p1;

assign r_V_146_fu_514_p1 = 44'd1601;

assign r_V_147_fu_508_p0 = sext_ln70_84_fu_33561_p1;

assign r_V_147_fu_508_p1 = 44'd1095;

assign r_V_148_fu_518_p0 = sext_ln70_81_fu_33548_p1;

assign r_V_148_fu_518_p1 = 49'd55758;

assign r_V_149_fu_493_p1 = 55'd7442488;

assign r_V_150_fu_531_p0 = sext_ln70_88_fu_34159_p1;

assign r_V_150_fu_531_p1 = 42'd495;

assign r_V_151_fu_517_p0 = sext_ln70_87_fu_34154_p1;

assign r_V_151_fu_517_p1 = 44'd17592186043304;

assign r_V_152_fu_516_p0 = sext_ln70_86_fu_34148_p1;

assign r_V_152_fu_516_p1 = 50'd97396;

assign r_V_153_fu_473_p0 = sext_ln70_86_fu_34148_p1;

assign r_V_153_fu_473_p1 = 50'd1125899906729295;

assign r_V_154_fu_523_p0 = sext_ln70_88_fu_34159_p1;

assign r_V_154_fu_523_p1 = 42'd372;

assign r_V_155_fu_483_p0 = sext_ln70_87_fu_34154_p1;

assign r_V_155_fu_483_p1 = 44'd17592186043249;

assign r_V_156_fu_34490_p2 = ($signed(sub_ln1273_10_fu_34473_p2) - $signed(sext_ln1273_21_fu_34486_p1));

assign r_V_157_fu_467_p0 = sext_ln70_86_fu_34148_p1;

assign r_V_157_fu_467_p1 = 50'd1125899906735636;

assign r_V_78_fu_527_p0 = sext_ln70_47_fu_17260_p1;

assign r_V_78_fu_527_p1 = 43'd8796093021384;

assign r_V_79_fu_484_p0 = sext_ln70_46_fu_17254_p1;

assign r_V_79_fu_484_p1 = 44'd17592186042992;

assign r_V_80_fu_509_p0 = sext_ln70_48_fu_17266_p1;

assign r_V_80_fu_509_p1 = 42'd427;

assign r_V_81_fu_489_p0 = sext_ln70_48_fu_17266_p1;

assign r_V_81_fu_489_p1 = 42'd482;

assign r_V_82_fu_497_p0 = sext_ln70_46_fu_17254_p1;

assign r_V_82_fu_497_p1 = 44'd17592186043065;

assign r_V_83_fu_507_p1 = 45'd2568;

assign r_V_84_fu_494_p1 = 40'd1099511627673;

assign r_V_85_fu_495_p0 = sext_ln70_47_fu_17260_p1;

assign r_V_85_fu_495_p1 = 43'd918;

assign r_V_86_fu_505_p1 = 45'd2170;

assign r_V_87_fu_538_p0 = sext_ln70_53_fu_17869_p1;

assign r_V_87_fu_538_p1 = 42'd410;

assign r_V_88_fu_498_p1 = 40'd1099511627665;

assign r_V_89_fu_482_p1 = 44'd17592186043166;

assign r_V_90_fu_480_p0 = sext_ln70_53_fu_17869_p1;

assign r_V_90_fu_480_p1 = 42'd4398046510682;

assign r_V_91_fu_18121_p2 = ($signed(sub_ln1273_fu_18103_p2) - $signed(sext_ln1273_13_fu_18117_p1));

assign r_V_92_fu_522_p0 = sext_ln70_53_fu_17869_p1;

assign r_V_92_fu_522_p1 = 42'd290;

assign r_V_93_fu_532_p1 = 43'd843;

assign r_V_94_fu_499_p1 = 39'd549755813843;

assign r_V_95_fu_503_p1 = 55'd36028797011701431;

assign r_V_96_fu_530_p1 = 44'd1428;

assign r_V_97_fu_504_p0 = sext_ln70_60_fu_18458_p1;

assign r_V_97_fu_504_p1 = 41'd135;

assign r_V_98_fu_501_p1 = 56'd14737058;

assign r_V_99_fu_465_p1 = 52'd4503599626520398;

assign r_V_fu_536_p0 = sext_ln70_48_fu_17266_p1;

assign r_V_fu_536_p1 = 42'd498;

assign ret_V_100_fu_29389_p2 = ($signed(sext_ln813_184_fu_29385_p1) + $signed(sext_ln813_183_fu_29382_p1));

assign ret_V_101_fu_29488_p2 = ($signed(sext_ln813_186_fu_29485_p1) + $signed(sext_ln813_185_fu_29482_p1));

assign ret_V_102_fu_29587_p2 = ($signed(sext_ln813_188_fu_29583_p1) + $signed(sext_ln813_187_fu_29580_p1));

assign ret_V_103_fu_29687_p2 = ($signed(sext_ln813_190_fu_29683_p1) + $signed(sext_ln813_189_fu_29680_p1));

assign ret_V_104_fu_29787_p2 = ($signed(sext_ln813_192_fu_29783_p1) + $signed(sext_ln813_191_fu_29780_p1));

assign ret_V_105_fu_29887_p2 = ($signed(sext_ln813_194_fu_29883_p1) + $signed(sext_ln813_193_fu_29880_p1));

assign ret_V_106_fu_29987_p2 = ($signed(sext_ln813_196_fu_29983_p1) + $signed(sext_ln813_195_fu_29980_p1));

assign ret_V_107_fu_30088_p2 = ($signed(sext_ln813_198_fu_30084_p1) + $signed(sext_ln813_197_fu_30080_p1));

assign ret_V_108_fu_30190_p2 = ($signed(sext_ln813_200_fu_30186_p1) + $signed(sext_ln813_199_fu_30182_p1));

assign ret_V_109_fu_30292_p2 = ($signed(sext_ln813_202_fu_30288_p1) + $signed(sext_ln813_201_fu_30284_p1));

assign ret_V_110_fu_30394_p2 = ($signed(sext_ln813_204_fu_30390_p1) + $signed(sext_ln813_203_fu_30386_p1));

assign ret_V_111_fu_30496_p2 = ($signed(sext_ln813_206_fu_30492_p1) + $signed(sext_ln813_205_fu_30488_p1));

assign ret_V_112_fu_30598_p2 = ($signed(sext_ln813_208_fu_30594_p1) + $signed(sext_ln813_207_fu_30590_p1));

assign ret_V_113_fu_30700_p2 = ($signed(sext_ln813_210_fu_30696_p1) + $signed(sext_ln813_209_fu_30692_p1));

assign ret_V_114_fu_30802_p2 = ($signed(sext_ln813_212_fu_30798_p1) + $signed(sext_ln813_211_fu_30794_p1));

assign ret_V_115_fu_30904_p2 = ($signed(sext_ln813_214_fu_30900_p1) + $signed(sext_ln813_213_fu_30896_p1));

assign ret_V_116_fu_31006_p2 = ($signed(sext_ln813_216_fu_31002_p1) + $signed(sext_ln813_215_fu_30998_p1));

assign ret_V_117_fu_31042_p2 = ($signed(sext_ln813_218_fu_31038_p1) + $signed(sext_ln813_217_fu_31034_p1));

assign ret_V_118_fu_31078_p2 = ($signed(sext_ln813_220_fu_31074_p1) + $signed(sext_ln813_219_fu_31070_p1));

assign ret_V_119_fu_31114_p2 = ($signed(sext_ln813_222_fu_31110_p1) + $signed(sext_ln813_221_fu_31106_p1));

assign ret_V_120_fu_31150_p2 = ($signed(sext_ln813_224_fu_31146_p1) + $signed(sext_ln813_223_fu_31142_p1));

assign ret_V_121_fu_31186_p2 = ($signed(sext_ln813_226_fu_31182_p1) + $signed(sext_ln813_225_fu_31178_p1));

assign ret_V_122_fu_31222_p2 = ($signed(sext_ln813_228_fu_31218_p1) + $signed(sext_ln813_227_fu_31214_p1));

assign ret_V_123_fu_31258_p2 = ($signed(sext_ln813_230_fu_31254_p1) + $signed(sext_ln813_229_fu_31250_p1));

assign ret_V_124_fu_31294_p2 = ($signed(sext_ln813_232_fu_31290_p1) + $signed(sext_ln813_231_fu_31286_p1));

assign ret_V_125_fu_35248_p2 = ($signed(sext_ln813_234_fu_35244_p1) + $signed(sext_ln813_233_fu_35240_p1));

assign ret_V_126_fu_35350_p2 = ($signed(sext_ln813_236_fu_35346_p1) + $signed(sext_ln813_235_fu_35342_p1));

assign ret_V_127_fu_35452_p2 = ($signed(sext_ln813_238_fu_35448_p1) + $signed(sext_ln813_237_fu_35444_p1));

assign ret_V_128_fu_35554_p2 = ($signed(sext_ln813_240_fu_35550_p1) + $signed(sext_ln813_239_fu_35546_p1));

assign ret_V_129_fu_35656_p2 = ($signed(sext_ln813_242_fu_35652_p1) + $signed(sext_ln813_241_fu_35648_p1));

assign ret_V_130_fu_35758_p2 = ($signed(sext_ln813_244_fu_35754_p1) + $signed(sext_ln813_243_fu_35750_p1));

assign ret_V_131_fu_35860_p2 = ($signed(sext_ln813_246_fu_35856_p1) + $signed(sext_ln813_245_fu_35852_p1));

assign ret_V_132_fu_35962_p2 = ($signed(sext_ln813_248_fu_35958_p1) + $signed(sext_ln813_247_fu_35954_p1));

assign ret_V_133_fu_36064_p2 = ($signed(sext_ln813_250_fu_36060_p1) + $signed(sext_ln813_249_fu_36056_p1));

assign ret_V_134_fu_36166_p2 = ($signed(sext_ln813_252_fu_36162_p1) + $signed(sext_ln813_251_fu_36158_p1));

assign ret_V_135_fu_36268_p2 = ($signed(sext_ln813_254_fu_36264_p1) + $signed(sext_ln813_253_fu_36260_p1));

assign ret_V_136_fu_36370_p2 = ($signed(sext_ln813_256_fu_36366_p1) + $signed(sext_ln813_255_fu_36362_p1));

assign ret_V_137_fu_36472_p2 = ($signed(sext_ln813_258_fu_36468_p1) + $signed(sext_ln813_257_fu_36464_p1));

assign ret_V_138_fu_36574_p2 = ($signed(sext_ln813_260_fu_36570_p1) + $signed(sext_ln813_259_fu_36566_p1));

assign ret_V_139_fu_36676_p2 = ($signed(sext_ln813_262_fu_36672_p1) + $signed(sext_ln813_261_fu_36668_p1));

assign ret_V_140_fu_36778_p2 = ($signed(sext_ln813_264_fu_36774_p1) + $signed(sext_ln813_263_fu_36770_p1));

assign ret_V_141_fu_36880_p2 = ($signed(sext_ln813_266_fu_36876_p1) + $signed(sext_ln813_265_fu_36872_p1));

assign ret_V_142_fu_36982_p2 = ($signed(sext_ln813_268_fu_36978_p1) + $signed(sext_ln813_267_fu_36974_p1));

assign ret_V_143_fu_39409_p2 = ($signed(sext_ln813_270_fu_39405_p1) + $signed(sext_ln813_269_fu_39402_p1));

assign ret_V_144_fu_39509_p2 = ($signed(sext_ln813_272_fu_39505_p1) + $signed(sext_ln813_271_fu_39502_p1));

assign ret_V_145_fu_39609_p2 = ($signed(sext_ln813_274_fu_39605_p1) + $signed(sext_ln813_273_fu_39602_p1));

assign ret_V_146_fu_39709_p2 = ($signed(sext_ln813_276_fu_39705_p1) + $signed(sext_ln813_275_fu_39702_p1));

assign ret_V_147_fu_39809_p2 = ($signed(sext_ln813_278_fu_39805_p1) + $signed(sext_ln813_277_fu_39802_p1));

assign ret_V_148_fu_39909_p2 = ($signed(sext_ln813_280_fu_39905_p1) + $signed(sext_ln813_279_fu_39902_p1));

assign ret_V_149_fu_40009_p2 = ($signed(sext_ln813_282_fu_40005_p1) + $signed(sext_ln813_281_fu_40002_p1));

assign ret_V_150_fu_40109_p2 = ($signed(sext_ln813_284_fu_40105_p1) + $signed(sext_ln813_283_fu_40102_p1));

assign ret_V_151_fu_40209_p2 = ($signed(sext_ln813_286_fu_40205_p1) + $signed(sext_ln813_285_fu_40202_p1));

assign ret_V_152_fu_40310_p2 = ($signed(sext_ln813_288_fu_40306_p1) + $signed(sext_ln813_287_fu_40302_p1));

assign ret_V_153_fu_40412_p2 = ($signed(sext_ln813_290_fu_40408_p1) + $signed(sext_ln813_289_fu_40404_p1));

assign ret_V_154_fu_40514_p2 = ($signed(sext_ln813_292_fu_40510_p1) + $signed(sext_ln813_291_fu_40506_p1));

assign ret_V_155_fu_40616_p2 = ($signed(sext_ln813_294_fu_40612_p1) + $signed(sext_ln813_293_fu_40608_p1));

assign ret_V_156_fu_40718_p2 = ($signed(sext_ln813_296_fu_40714_p1) + $signed(sext_ln813_295_fu_40710_p1));

assign ret_V_157_fu_40820_p2 = ($signed(sext_ln813_298_fu_40816_p1) + $signed(sext_ln813_297_fu_40812_p1));

assign ret_V_158_fu_40922_p2 = ($signed(sext_ln813_300_fu_40918_p1) + $signed(sext_ln813_299_fu_40914_p1));

assign ret_V_159_fu_41024_p2 = ($signed(sext_ln813_302_fu_41020_p1) + $signed(sext_ln813_301_fu_41016_p1));

assign ret_V_160_fu_41126_p2 = ($signed(sext_ln813_304_fu_41122_p1) + $signed(sext_ln813_303_fu_41118_p1));

assign ret_V_81_fu_23724_p2 = ($signed(sext_ln813_153_fu_23720_p1) + $signed(33'd8589885299));

assign ret_V_82_fu_23822_p2 = ($signed(sext_ln813_154_fu_23818_p1) + $signed(33'd8589341049));

assign ret_V_83_fu_23920_p2 = ($signed(sext_ln813_155_fu_23916_p1) + $signed(33'd8589929421));

assign ret_V_84_fu_24018_p2 = ($signed(sext_ln813_156_fu_24014_p1) + $signed(33'd6442053));

assign ret_V_85_fu_24116_p2 = ($signed(sext_ln813_157_fu_24112_p1) + $signed(33'd8589930485));

assign ret_V_86_fu_24214_p2 = ($signed(sext_ln813_158_fu_24210_p1) + $signed(33'd8589779773));

assign ret_V_87_fu_24312_p2 = ($signed(sext_ln813_159_fu_24308_p1) + $signed(33'd8589720800));

assign ret_V_88_fu_24410_p2 = ($signed(sext_ln813_160_fu_24406_p1) + $signed(33'd19328802));

assign ret_V_89_fu_24512_p2 = ($signed(sext_ln813_162_fu_24508_p1) + $signed(sext_ln813_161_fu_24504_p1));

assign ret_V_90_fu_24614_p2 = ($signed(sext_ln813_164_fu_24610_p1) + $signed(sext_ln813_163_fu_24606_p1));

assign ret_V_91_fu_24716_p2 = ($signed(sext_ln813_166_fu_24712_p1) + $signed(sext_ln813_165_fu_24708_p1));

assign ret_V_92_fu_24818_p2 = ($signed(sext_ln813_168_fu_24814_p1) + $signed(sext_ln813_167_fu_24810_p1));

assign ret_V_93_fu_24920_p2 = ($signed(sext_ln813_170_fu_24916_p1) + $signed(sext_ln813_169_fu_24912_p1));

assign ret_V_94_fu_25022_p2 = ($signed(sext_ln813_172_fu_25018_p1) + $signed(sext_ln813_171_fu_25014_p1));

assign ret_V_95_fu_25124_p2 = ($signed(sext_ln813_174_fu_25120_p1) + $signed(sext_ln813_173_fu_25116_p1));

assign ret_V_96_fu_25226_p2 = ($signed(sext_ln813_176_fu_25222_p1) + $signed(sext_ln813_175_fu_25218_p1));

assign ret_V_97_fu_25328_p2 = ($signed(sext_ln813_178_fu_25324_p1) + $signed(sext_ln813_177_fu_25320_p1));

assign ret_V_98_fu_29190_p2 = ($signed(sext_ln813_180_fu_29187_p1) + $signed(sext_ln813_179_fu_29184_p1));

assign ret_V_99_fu_29289_p2 = ($signed(sext_ln813_182_fu_29285_p1) + $signed(sext_ln813_181_fu_29282_p1));

assign ret_V_fu_23626_p2 = ($signed(sext_ln813_fu_23622_p1) + $signed(33'd5264183));

assign rhs_100_fu_25449_p3 = ((or_ln346_100_reg_42166[0:0] == 1'b1) ? select_ln346_182_fu_25442_p3 : sext_ln856_96_fu_25439_p1);

assign rhs_101_fu_21836_p3 = ((or_ln346_101_fu_21830_p2[0:0] == 1'b1) ? select_ln346_183_fu_21822_p3 : p_Val2_466_fu_21706_p2);

assign rhs_102_fu_25466_p3 = ((or_ln346_102_reg_42187[0:0] == 1'b1) ? select_ln346_184_fu_25459_p3 : sext_ln856_97_fu_25456_p1);

assign rhs_103_fu_25483_p3 = ((or_ln346_103_reg_42202[0:0] == 1'b1) ? select_ln346_185_fu_25476_p3 : sext_ln856_98_fu_25473_p1);

assign rhs_104_fu_25500_p3 = ((or_ln346_104_reg_42217[0:0] == 1'b1) ? select_ln346_186_fu_25493_p3 : sext_ln856_99_fu_25490_p1);

assign rhs_105_fu_25517_p3 = ((or_ln346_105_reg_42232[0:0] == 1'b1) ? select_ln346_187_fu_25510_p3 : sext_ln856_100_fu_25507_p1);

assign rhs_106_fu_25534_p3 = ((or_ln346_106_reg_42247[0:0] == 1'b1) ? select_ln346_188_fu_25527_p3 : sext_ln856_101_fu_25524_p1);

assign rhs_107_fu_25658_p3 = ((or_ln346_107_fu_25652_p2[0:0] == 1'b1) ? select_ln346_189_fu_25644_p3 : sext_ln856_102_fu_25541_p1);

assign rhs_108_fu_25783_p3 = ((or_ln346_108_fu_25777_p2[0:0] == 1'b1) ? select_ln346_190_fu_25769_p3 : sext_ln856_103_fu_25666_p1);

assign rhs_109_fu_25908_p3 = ((or_ln346_109_fu_25902_p2[0:0] == 1'b1) ? select_ln346_191_fu_25894_p3 : sext_ln856_104_fu_25791_p1);

assign rhs_110_fu_26033_p3 = ((or_ln346_110_fu_26027_p2[0:0] == 1'b1) ? select_ln346_192_fu_26019_p3 : sext_ln856_105_fu_25916_p1);

assign rhs_111_fu_26158_p3 = ((or_ln346_111_fu_26152_p2[0:0] == 1'b1) ? select_ln346_193_fu_26144_p3 : sext_ln856_106_fu_26041_p1);

assign rhs_112_fu_26283_p3 = ((or_ln346_112_fu_26277_p2[0:0] == 1'b1) ? select_ln346_194_fu_26269_p3 : sext_ln856_107_fu_26166_p1);

assign rhs_113_fu_26301_p3 = ((or_ln346_113_reg_42448[0:0] == 1'b1) ? select_ln346_195_fu_26294_p3 : sext_ln856_108_fu_26291_p1);

assign rhs_114_fu_26425_p3 = ((or_ln346_114_fu_26419_p2[0:0] == 1'b1) ? select_ln346_196_fu_26411_p3 : sext_ln856_109_fu_26308_p1);

assign rhs_115_fu_26550_p3 = ((or_ln346_115_fu_26544_p2[0:0] == 1'b1) ? select_ln346_197_fu_26536_p3 : sext_ln856_110_fu_26433_p1);

assign rhs_116_fu_26695_p3 = ((or_ln346_116_fu_26689_p2[0:0] == 1'b1) ? select_ln346_198_fu_26681_p3 : p_Val2_511_fu_26564_p2);

assign rhs_117_fu_26844_p3 = ((or_ln346_117_fu_26838_p2[0:0] == 1'b1) ? select_ln346_199_fu_26830_p3 : sext_ln856_111_fu_26715_p1);

assign rhs_118_fu_26993_p3 = ((or_ln346_118_fu_26987_p2[0:0] == 1'b1) ? select_ln346_200_fu_26979_p3 : sext_ln856_112_fu_26864_p1);

assign rhs_119_fu_27142_p3 = ((or_ln346_119_fu_27136_p2[0:0] == 1'b1) ? select_ln346_201_fu_27128_p3 : sext_ln856_113_fu_27013_p1);

assign rhs_120_fu_27291_p3 = ((or_ln346_120_fu_27285_p2[0:0] == 1'b1) ? select_ln346_202_fu_27277_p3 : sext_ln856_114_fu_27162_p1);

assign rhs_121_fu_27440_p3 = ((or_ln346_121_fu_27434_p2[0:0] == 1'b1) ? select_ln346_203_fu_27426_p3 : sext_ln856_115_fu_27311_p1);

assign rhs_122_fu_27589_p3 = ((or_ln346_122_fu_27583_p2[0:0] == 1'b1) ? select_ln346_204_fu_27575_p3 : sext_ln856_116_fu_27460_p1);

assign rhs_123_fu_27738_p3 = ((or_ln346_123_fu_27732_p2[0:0] == 1'b1) ? select_ln346_205_fu_27724_p3 : sext_ln856_117_fu_27609_p1);

assign rhs_124_fu_27887_p3 = ((or_ln346_124_fu_27881_p2[0:0] == 1'b1) ? select_ln346_206_fu_27873_p3 : sext_ln856_118_fu_27758_p1);

assign rhs_125_fu_31332_p3 = ((or_ln346_125_reg_42840[0:0] == 1'b1) ? select_ln346_207_fu_31325_p3 : sext_ln856_119_fu_31322_p1);

assign rhs_126_fu_31456_p3 = ((or_ln346_126_fu_31450_p2[0:0] == 1'b1) ? select_ln346_208_fu_31442_p3 : sext_ln856_120_fu_31339_p1);

assign rhs_127_fu_31581_p3 = ((or_ln346_127_fu_31575_p2[0:0] == 1'b1) ? select_ln346_209_fu_31567_p3 : sext_ln856_121_fu_31464_p1);

assign rhs_128_fu_31706_p3 = ((or_ln346_128_fu_31700_p2[0:0] == 1'b1) ? select_ln346_210_fu_31692_p3 : sext_ln856_122_fu_31589_p1);

assign rhs_129_fu_31831_p3 = ((or_ln346_129_fu_31825_p2[0:0] == 1'b1) ? select_ln346_211_fu_31817_p3 : sext_ln856_123_fu_31714_p1);

assign rhs_130_fu_31956_p3 = ((or_ln346_130_fu_31950_p2[0:0] == 1'b1) ? select_ln346_212_fu_31942_p3 : sext_ln856_124_fu_31839_p1);

assign rhs_131_fu_32081_p3 = ((or_ln346_131_fu_32075_p2[0:0] == 1'b1) ? select_ln346_213_fu_32067_p3 : sext_ln856_125_fu_31964_p1);

assign rhs_132_fu_32206_p3 = ((or_ln346_132_fu_32200_p2[0:0] == 1'b1) ? select_ln346_214_fu_32192_p3 : sext_ln856_126_fu_32089_p1);

assign rhs_133_fu_32331_p3 = ((or_ln346_133_fu_32325_p2[0:0] == 1'b1) ? select_ln346_215_fu_32317_p3 : sext_ln856_127_fu_32214_p1);

assign rhs_134_fu_32480_p3 = ((or_ln346_134_fu_32474_p2[0:0] == 1'b1) ? select_ln346_216_fu_32466_p3 : sext_ln856_128_fu_32351_p1);

assign rhs_135_fu_32629_p3 = ((or_ln346_135_fu_32623_p2[0:0] == 1'b1) ? select_ln346_217_fu_32615_p3 : sext_ln856_129_fu_32500_p1);

assign rhs_136_fu_32778_p3 = ((or_ln346_136_fu_32772_p2[0:0] == 1'b1) ? select_ln346_218_fu_32764_p3 : sext_ln856_130_fu_32649_p1);

assign rhs_137_fu_32927_p3 = ((or_ln346_137_fu_32921_p2[0:0] == 1'b1) ? select_ln346_219_fu_32913_p3 : sext_ln856_131_fu_32798_p1);

assign rhs_138_fu_33076_p3 = ((or_ln346_138_fu_33070_p2[0:0] == 1'b1) ? select_ln346_220_fu_33062_p3 : sext_ln856_132_fu_32947_p1);

assign rhs_139_fu_33225_p3 = ((or_ln346_139_fu_33219_p2[0:0] == 1'b1) ? select_ln346_221_fu_33211_p3 : sext_ln856_133_fu_33096_p1);

assign rhs_140_fu_33374_p3 = ((or_ln346_140_fu_33368_p2[0:0] == 1'b1) ? select_ln346_222_fu_33360_p3 : sext_ln856_134_fu_33245_p1);

assign rhs_141_fu_33523_p3 = ((or_ln346_141_fu_33517_p2[0:0] == 1'b1) ? select_ln346_223_fu_33509_p3 : sext_ln856_135_fu_33394_p1);

assign rhs_142_fu_33541_p3 = ((or_ln346_142_reg_43335[0:0] == 1'b1) ? select_ln346_224_fu_33534_p3 : sext_ln856_136_fu_33531_p1);

assign rhs_143_fu_37190_p3 = ((or_ln346_143_fu_37184_p2[0:0] == 1'b1) ? select_ln346_225_fu_37176_p3 : p_Val2_592_reg_43532);

assign rhs_144_fu_37314_p3 = ((or_ln346_144_fu_37308_p2[0:0] == 1'b1) ? select_ln346_226_fu_37300_p3 : sext_ln856_137_fu_37197_p1);

assign rhs_145_fu_37439_p3 = ((or_ln346_145_fu_37433_p2[0:0] == 1'b1) ? select_ln346_227_fu_37425_p3 : sext_ln856_138_fu_37322_p1);

assign rhs_146_fu_37564_p3 = ((or_ln346_146_fu_37558_p2[0:0] == 1'b1) ? select_ln346_228_fu_37550_p3 : sext_ln856_139_fu_37447_p1);

assign rhs_147_fu_37689_p3 = ((or_ln346_147_fu_37683_p2[0:0] == 1'b1) ? select_ln346_229_fu_37675_p3 : sext_ln856_140_fu_37572_p1);

assign rhs_148_fu_37814_p3 = ((or_ln346_148_fu_37808_p2[0:0] == 1'b1) ? select_ln346_230_fu_37800_p3 : sext_ln856_141_fu_37697_p1);

assign rhs_149_fu_37939_p3 = ((or_ln346_149_fu_37933_p2[0:0] == 1'b1) ? select_ln346_231_fu_37925_p3 : sext_ln856_142_fu_37822_p1);

assign rhs_150_fu_38064_p3 = ((or_ln346_150_fu_38058_p2[0:0] == 1'b1) ? select_ln346_232_fu_38050_p3 : sext_ln856_143_fu_37947_p1);

assign rhs_151_fu_38189_p3 = ((or_ln346_151_fu_38183_p2[0:0] == 1'b1) ? select_ln346_233_fu_38175_p3 : sext_ln856_144_fu_38072_p1);

assign rhs_152_fu_38334_p3 = ((or_ln346_152_fu_38328_p2[0:0] == 1'b1) ? select_ln346_234_fu_38320_p3 : p_Val2_619_fu_38203_p2);

assign rhs_153_fu_38483_p3 = ((or_ln346_153_fu_38477_p2[0:0] == 1'b1) ? select_ln346_235_fu_38469_p3 : sext_ln856_145_fu_38354_p1);

assign rhs_154_fu_38632_p3 = ((or_ln346_154_fu_38626_p2[0:0] == 1'b1) ? select_ln346_236_fu_38618_p3 : sext_ln856_146_fu_38503_p1);

assign rhs_155_fu_38781_p3 = ((or_ln346_155_fu_38775_p2[0:0] == 1'b1) ? select_ln346_237_fu_38767_p3 : sext_ln856_147_fu_38652_p1);

assign rhs_156_fu_38930_p3 = ((or_ln346_156_fu_38924_p2[0:0] == 1'b1) ? select_ln346_238_fu_38916_p3 : sext_ln856_148_fu_38801_p1);

assign rhs_157_fu_39079_p3 = ((or_ln346_157_fu_39073_p2[0:0] == 1'b1) ? select_ln346_239_fu_39065_p3 : sext_ln856_149_fu_38950_p1);

assign rhs_158_fu_39228_p3 = ((or_ln346_158_fu_39222_p2[0:0] == 1'b1) ? select_ln346_240_fu_39214_p3 : sext_ln856_150_fu_39099_p1);

assign rhs_159_fu_39246_p3 = ((or_ln346_159_reg_44012[0:0] == 1'b1) ? select_ln346_241_fu_39239_p3 : sext_ln856_151_fu_39236_p1);

assign rhs_160_fu_39394_p3 = ((or_ln346_160_fu_39388_p2[0:0] == 1'b1) ? select_ln346_242_fu_39380_p3 : sext_ln856_152_fu_39265_p1);

assign rhs_81_fu_19208_p3 = ((or_ln346_81_fu_19202_p2[0:0] == 1'b1) ? select_ln346_163_fu_19194_p3 : sext_ln856_78_fu_19091_p1);

assign rhs_82_fu_19333_p3 = ((or_ln346_82_fu_19327_p2[0:0] == 1'b1) ? select_ln346_164_fu_19319_p3 : sext_ln856_79_fu_19216_p1);

assign rhs_83_fu_19458_p3 = ((or_ln346_83_fu_19452_p2[0:0] == 1'b1) ? select_ln346_165_fu_19444_p3 : sext_ln856_80_fu_19341_p1);

assign rhs_84_fu_19583_p3 = ((or_ln346_84_fu_19577_p2[0:0] == 1'b1) ? select_ln346_166_fu_19569_p3 : sext_ln856_81_fu_19466_p1);

assign rhs_85_fu_19708_p3 = ((or_ln346_85_fu_19702_p2[0:0] == 1'b1) ? select_ln346_167_fu_19694_p3 : sext_ln856_82_fu_19591_p1);

assign rhs_86_fu_19833_p3 = ((or_ln346_86_fu_19827_p2[0:0] == 1'b1) ? select_ln346_168_fu_19819_p3 : sext_ln856_83_fu_19716_p1);

assign rhs_87_fu_19958_p3 = ((or_ln346_87_fu_19952_p2[0:0] == 1'b1) ? select_ln346_169_fu_19944_p3 : sext_ln856_84_fu_19841_p1);

assign rhs_88_fu_20083_p3 = ((or_ln346_88_fu_20077_p2[0:0] == 1'b1) ? select_ln346_170_fu_20069_p3 : sext_ln856_85_fu_19966_p1);

assign rhs_89_fu_20232_p3 = ((or_ln346_89_fu_20226_p2[0:0] == 1'b1) ? select_ln346_171_fu_20218_p3 : sext_ln856_86_fu_20103_p1);

assign rhs_90_fu_20381_p3 = ((or_ln346_90_fu_20375_p2[0:0] == 1'b1) ? select_ln346_172_fu_20367_p3 : sext_ln856_87_fu_20252_p1);

assign rhs_91_fu_20530_p3 = ((or_ln346_91_fu_20524_p2[0:0] == 1'b1) ? select_ln346_173_fu_20516_p3 : sext_ln856_88_fu_20401_p1);

assign rhs_92_fu_20679_p3 = ((or_ln346_92_fu_20673_p2[0:0] == 1'b1) ? select_ln346_174_fu_20665_p3 : sext_ln856_89_fu_20550_p1);

assign rhs_93_fu_20828_p3 = ((or_ln346_93_fu_20822_p2[0:0] == 1'b1) ? select_ln346_175_fu_20814_p3 : sext_ln856_90_fu_20699_p1);

assign rhs_94_fu_20846_p3 = ((or_ln346_94_reg_41767[0:0] == 1'b1) ? select_ln346_176_fu_20839_p3 : sext_ln856_91_fu_20836_p1);

assign rhs_95_fu_20994_p3 = ((or_ln346_95_fu_20988_p2[0:0] == 1'b1) ? select_ln346_177_fu_20980_p3 : sext_ln856_92_fu_20865_p1);

assign rhs_96_fu_21143_p3 = ((or_ln346_96_fu_21137_p2[0:0] == 1'b1) ? select_ln346_178_fu_21129_p3 : sext_ln856_93_fu_21014_p1);

assign rhs_97_fu_21292_p3 = ((or_ln346_97_fu_21286_p2[0:0] == 1'b1) ? select_ln346_179_fu_21278_p3 : sext_ln856_94_fu_21163_p1);

assign rhs_98_fu_21437_p3 = ((or_ln346_98_fu_21431_p2[0:0] == 1'b1) ? select_ln346_180_fu_21423_p3 : p_Val2_457_fu_21306_p2);

assign rhs_99_fu_25432_p3 = ((or_ln346_99_reg_42151[0:0] == 1'b1) ? select_ln346_181_fu_25425_p3 : sext_ln856_95_fu_25422_p1);

assign rhs_fu_19083_p3 = ((or_ln346_fu_19077_p2[0:0] == 1'b1) ? select_ln346_fu_19069_p3 : sext_ln856_fu_18966_p1);

assign select_ln302_163_fu_23794_p3 = ((xor_ln302_163_fu_23776_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_647_fu_23738_p2);

assign select_ln302_165_fu_23892_p3 = ((xor_ln302_165_fu_23874_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_649_fu_23836_p2);

assign select_ln302_167_fu_23990_p3 = ((xor_ln302_167_fu_23972_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_651_fu_23934_p2);

assign select_ln302_169_fu_24088_p3 = ((xor_ln302_169_fu_24070_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_653_fu_24032_p2);

assign select_ln302_171_fu_24186_p3 = ((xor_ln302_171_fu_24168_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_655_fu_24130_p2);

assign select_ln302_173_fu_24284_p3 = ((xor_ln302_173_fu_24266_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_657_fu_24228_p2);

assign select_ln302_175_fu_24382_p3 = ((xor_ln302_175_fu_24364_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_659_fu_24326_p2);

assign select_ln302_177_fu_24480_p3 = ((xor_ln302_177_fu_24462_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_661_fu_24424_p2);

assign select_ln302_179_fu_24582_p3 = ((xor_ln302_179_fu_24564_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_663_fu_24526_p2);

assign select_ln302_181_fu_24684_p3 = ((xor_ln302_181_fu_24666_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_665_fu_24628_p2);

assign select_ln302_183_fu_24786_p3 = ((xor_ln302_183_fu_24768_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_667_fu_24730_p2);

assign select_ln302_185_fu_24888_p3 = ((xor_ln302_185_fu_24870_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_669_fu_24832_p2);

assign select_ln302_187_fu_24990_p3 = ((xor_ln302_187_fu_24972_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_671_fu_24934_p2);

assign select_ln302_189_fu_25092_p3 = ((xor_ln302_189_fu_25074_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_673_fu_25036_p2);

assign select_ln302_191_fu_25194_p3 = ((xor_ln302_191_fu_25176_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_675_fu_25138_p2);

assign select_ln302_193_fu_25296_p3 = ((xor_ln302_193_fu_25278_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_677_fu_25240_p2);

assign select_ln302_195_fu_25398_p3 = ((xor_ln302_195_fu_25380_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_679_fu_25342_p2);

assign select_ln302_197_fu_29258_p3 = ((xor_ln302_197_fu_29240_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_681_fu_29204_p2);

assign select_ln302_199_fu_29358_p3 = ((xor_ln302_199_fu_29340_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_683_fu_29303_p2);

assign select_ln302_201_fu_29458_p3 = ((xor_ln302_201_fu_29440_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_685_fu_29403_p2);

assign select_ln302_203_fu_29556_p3 = ((xor_ln302_203_fu_29538_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_687_fu_29502_p2);

assign select_ln302_205_fu_29656_p3 = ((xor_ln302_205_fu_29638_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_689_fu_29601_p2);

assign select_ln302_207_fu_29756_p3 = ((xor_ln302_207_fu_29738_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_691_fu_29701_p2);

assign select_ln302_209_fu_29856_p3 = ((xor_ln302_209_fu_29838_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_693_fu_29801_p2);

assign select_ln302_211_fu_29956_p3 = ((xor_ln302_211_fu_29938_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_695_fu_29901_p2);

assign select_ln302_213_fu_30056_p3 = ((xor_ln302_213_fu_30038_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_697_fu_30001_p2);

assign select_ln302_215_fu_30158_p3 = ((xor_ln302_215_fu_30140_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_699_fu_30102_p2);

assign select_ln302_217_fu_30260_p3 = ((xor_ln302_217_fu_30242_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_701_fu_30204_p2);

assign select_ln302_219_fu_30362_p3 = ((xor_ln302_219_fu_30344_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_703_fu_30306_p2);

assign select_ln302_221_fu_30464_p3 = ((xor_ln302_221_fu_30446_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_705_fu_30408_p2);

assign select_ln302_223_fu_30566_p3 = ((xor_ln302_223_fu_30548_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_707_fu_30510_p2);

assign select_ln302_225_fu_30668_p3 = ((xor_ln302_225_fu_30650_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_709_fu_30612_p2);

assign select_ln302_227_fu_30770_p3 = ((xor_ln302_227_fu_30752_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_711_fu_30714_p2);

assign select_ln302_229_fu_30872_p3 = ((xor_ln302_229_fu_30854_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_713_fu_30816_p2);

assign select_ln302_231_fu_30974_p3 = ((xor_ln302_231_fu_30956_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_715_fu_30918_p2);

assign select_ln302_233_fu_34754_p3 = ((xor_ln302_233_fu_34738_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_717_reg_43347);

assign select_ln302_235_fu_34812_p3 = ((xor_ln302_235_fu_34796_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_719_reg_43367);

assign select_ln302_237_fu_34870_p3 = ((xor_ln302_237_fu_34854_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_721_reg_43387);

assign select_ln302_239_fu_34928_p3 = ((xor_ln302_239_fu_34912_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_723_reg_43407);

assign select_ln302_241_fu_34986_p3 = ((xor_ln302_241_fu_34970_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_725_reg_43427);

assign select_ln302_243_fu_35044_p3 = ((xor_ln302_243_fu_35028_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_727_reg_43447);

assign select_ln302_245_fu_35102_p3 = ((xor_ln302_245_fu_35086_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_729_reg_43467);

assign select_ln302_247_fu_35160_p3 = ((xor_ln302_247_fu_35144_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_731_reg_43487);

assign select_ln302_249_fu_35218_p3 = ((xor_ln302_249_fu_35202_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_733_reg_43507);

assign select_ln302_251_fu_35318_p3 = ((xor_ln302_251_fu_35300_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_735_fu_35262_p2);

assign select_ln302_253_fu_35420_p3 = ((xor_ln302_253_fu_35402_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_737_fu_35364_p2);

assign select_ln302_255_fu_35522_p3 = ((xor_ln302_255_fu_35504_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_739_fu_35466_p2);

assign select_ln302_257_fu_35624_p3 = ((xor_ln302_257_fu_35606_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_741_fu_35568_p2);

assign select_ln302_259_fu_35726_p3 = ((xor_ln302_259_fu_35708_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_743_fu_35670_p2);

assign select_ln302_261_fu_35828_p3 = ((xor_ln302_261_fu_35810_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_745_fu_35772_p2);

assign select_ln302_263_fu_35930_p3 = ((xor_ln302_263_fu_35912_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_747_fu_35874_p2);

assign select_ln302_265_fu_36032_p3 = ((xor_ln302_265_fu_36014_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_749_fu_35976_p2);

assign select_ln302_267_fu_36134_p3 = ((xor_ln302_267_fu_36116_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_751_fu_36078_p2);

assign select_ln302_269_fu_36236_p3 = ((xor_ln302_269_fu_36218_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_753_fu_36180_p2);

assign select_ln302_271_fu_36338_p3 = ((xor_ln302_271_fu_36320_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_755_fu_36282_p2);

assign select_ln302_273_fu_36440_p3 = ((xor_ln302_273_fu_36422_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_757_fu_36384_p2);

assign select_ln302_275_fu_36542_p3 = ((xor_ln302_275_fu_36524_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_759_fu_36486_p2);

assign select_ln302_277_fu_36644_p3 = ((xor_ln302_277_fu_36626_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_761_fu_36588_p2);

assign select_ln302_279_fu_36746_p3 = ((xor_ln302_279_fu_36728_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_763_fu_36690_p2);

assign select_ln302_281_fu_36848_p3 = ((xor_ln302_281_fu_36830_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_765_fu_36792_p2);

assign select_ln302_283_fu_36950_p3 = ((xor_ln302_283_fu_36932_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_767_fu_36894_p2);

assign select_ln302_285_fu_37052_p3 = ((xor_ln302_285_fu_37034_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_769_fu_36996_p2);

assign select_ln302_287_fu_39478_p3 = ((xor_ln302_287_fu_39460_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_771_fu_39423_p2);

assign select_ln302_289_fu_39578_p3 = ((xor_ln302_289_fu_39560_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_773_fu_39523_p2);

assign select_ln302_291_fu_39678_p3 = ((xor_ln302_291_fu_39660_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_775_fu_39623_p2);

assign select_ln302_293_fu_39778_p3 = ((xor_ln302_293_fu_39760_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_777_fu_39723_p2);

assign select_ln302_295_fu_39878_p3 = ((xor_ln302_295_fu_39860_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_779_fu_39823_p2);

assign select_ln302_297_fu_39978_p3 = ((xor_ln302_297_fu_39960_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_781_fu_39923_p2);

assign select_ln302_299_fu_40078_p3 = ((xor_ln302_299_fu_40060_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_783_fu_40023_p2);

assign select_ln302_301_fu_40178_p3 = ((xor_ln302_301_fu_40160_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_785_fu_40123_p2);

assign select_ln302_303_fu_40278_p3 = ((xor_ln302_303_fu_40260_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_787_fu_40223_p2);

assign select_ln302_305_fu_40380_p3 = ((xor_ln302_305_fu_40362_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_789_fu_40324_p2);

assign select_ln302_306_fu_40396_p3 = ((or_ln302_152_fu_40374_p2[0:0] == 1'b1) ? select_ln302_305_fu_40380_p3 : select_ln350_152_fu_40388_p3);

assign select_ln302_307_fu_40482_p3 = ((xor_ln302_307_fu_40464_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_791_fu_40426_p2);

assign select_ln302_308_fu_40498_p3 = ((or_ln302_153_fu_40476_p2[0:0] == 1'b1) ? select_ln302_307_fu_40482_p3 : select_ln350_153_fu_40490_p3);

assign select_ln302_309_fu_40584_p3 = ((xor_ln302_309_fu_40566_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_793_fu_40528_p2);

assign select_ln302_310_fu_40600_p3 = ((or_ln302_154_fu_40578_p2[0:0] == 1'b1) ? select_ln302_309_fu_40584_p3 : select_ln350_154_fu_40592_p3);

assign select_ln302_311_fu_40686_p3 = ((xor_ln302_311_fu_40668_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_795_fu_40630_p2);

assign select_ln302_312_fu_40702_p3 = ((or_ln302_155_fu_40680_p2[0:0] == 1'b1) ? select_ln302_311_fu_40686_p3 : select_ln350_155_fu_40694_p3);

assign select_ln302_313_fu_40788_p3 = ((xor_ln302_313_fu_40770_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_797_fu_40732_p2);

assign select_ln302_314_fu_40804_p3 = ((or_ln302_156_fu_40782_p2[0:0] == 1'b1) ? select_ln302_313_fu_40788_p3 : select_ln350_156_fu_40796_p3);

assign select_ln302_315_fu_40890_p3 = ((xor_ln302_315_fu_40872_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_799_fu_40834_p2);

assign select_ln302_316_fu_40906_p3 = ((or_ln302_157_fu_40884_p2[0:0] == 1'b1) ? select_ln302_315_fu_40890_p3 : select_ln350_157_fu_40898_p3);

assign select_ln302_317_fu_40992_p3 = ((xor_ln302_317_fu_40974_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_801_fu_40936_p2);

assign select_ln302_318_fu_41008_p3 = ((or_ln302_158_fu_40986_p2[0:0] == 1'b1) ? select_ln302_317_fu_40992_p3 : select_ln350_158_fu_41000_p3);

assign select_ln302_319_fu_41094_p3 = ((xor_ln302_319_fu_41076_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_803_fu_41038_p2);

assign select_ln302_320_fu_41110_p3 = ((or_ln302_159_fu_41088_p2[0:0] == 1'b1) ? select_ln302_319_fu_41094_p3 : select_ln350_159_fu_41102_p3);

assign select_ln302_321_fu_41196_p3 = ((xor_ln302_321_fu_41178_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_805_fu_41140_p2);

assign select_ln302_322_fu_41212_p3 = ((or_ln302_160_fu_41190_p2[0:0] == 1'b1) ? select_ln302_321_fu_41196_p3 : select_ln350_160_fu_41204_p3);

assign select_ln302_fu_23696_p3 = ((xor_ln302_fu_23678_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_645_fu_23640_p2);

assign select_ln346_163_fu_19194_p3 = ((overflow_162_fu_19165_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_164_fu_19319_p3 = ((overflow_163_fu_19290_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_165_fu_19444_p3 = ((overflow_164_fu_19415_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_166_fu_19569_p3 = ((overflow_165_fu_19540_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_167_fu_19694_p3 = ((overflow_166_fu_19665_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_168_fu_19819_p3 = ((overflow_167_fu_19790_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_169_fu_19944_p3 = ((overflow_168_fu_19915_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_170_fu_20069_p3 = ((overflow_169_fu_20040_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_171_fu_20218_p3 = ((overflow_170_fu_20189_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_172_fu_20367_p3 = ((overflow_171_fu_20338_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_173_fu_20516_p3 = ((overflow_172_fu_20487_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_174_fu_20665_p3 = ((overflow_173_fu_20636_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_175_fu_20814_p3 = ((overflow_174_fu_20785_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_176_fu_20839_p3 = ((overflow_175_reg_41762[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_177_fu_20980_p3 = ((overflow_176_fu_20951_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_178_fu_21129_p3 = ((overflow_177_fu_21100_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_179_fu_21278_p3 = ((overflow_178_fu_21249_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_180_fu_21423_p3 = ((overflow_179_fu_21394_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_181_fu_25425_p3 = ((overflow_180_reg_42146[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_182_fu_25442_p3 = ((overflow_181_reg_42161[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_183_fu_21822_p3 = ((overflow_182_fu_21793_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_184_fu_25459_p3 = ((overflow_183_reg_42182[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_185_fu_25476_p3 = ((overflow_184_reg_42197[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_186_fu_25493_p3 = ((overflow_185_reg_42212[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_187_fu_25510_p3 = ((overflow_186_reg_42227[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_188_fu_25527_p3 = ((overflow_187_reg_42242[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_189_fu_25644_p3 = ((overflow_188_fu_25615_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_190_fu_25769_p3 = ((overflow_189_fu_25740_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_191_fu_25894_p3 = ((overflow_190_fu_25865_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_192_fu_26019_p3 = ((overflow_191_fu_25990_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_193_fu_26144_p3 = ((overflow_192_fu_26115_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_194_fu_26269_p3 = ((overflow_193_fu_26240_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_195_fu_26294_p3 = ((overflow_194_reg_42443[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_196_fu_26411_p3 = ((overflow_195_fu_26382_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_197_fu_26536_p3 = ((overflow_196_fu_26507_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_198_fu_26681_p3 = ((overflow_197_fu_26652_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_199_fu_26830_p3 = ((overflow_198_fu_26801_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_200_fu_26979_p3 = ((overflow_199_fu_26950_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_201_fu_27128_p3 = ((overflow_200_fu_27099_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_202_fu_27277_p3 = ((overflow_201_fu_27248_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_203_fu_27426_p3 = ((overflow_202_fu_27397_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_204_fu_27575_p3 = ((overflow_203_fu_27546_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_205_fu_27724_p3 = ((overflow_204_fu_27695_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_206_fu_27873_p3 = ((overflow_205_fu_27844_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_207_fu_31325_p3 = ((overflow_206_reg_42835[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_208_fu_31442_p3 = ((overflow_207_fu_31413_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_209_fu_31567_p3 = ((overflow_208_fu_31538_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_210_fu_31692_p3 = ((overflow_209_fu_31663_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_211_fu_31817_p3 = ((overflow_210_fu_31788_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_212_fu_31942_p3 = ((overflow_211_fu_31913_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_213_fu_32067_p3 = ((overflow_212_fu_32038_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_214_fu_32192_p3 = ((overflow_213_fu_32163_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_215_fu_32317_p3 = ((overflow_214_fu_32288_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_216_fu_32466_p3 = ((overflow_215_fu_32437_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_217_fu_32615_p3 = ((overflow_216_fu_32586_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_218_fu_32764_p3 = ((overflow_217_fu_32735_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_219_fu_32913_p3 = ((overflow_218_fu_32884_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_220_fu_33062_p3 = ((overflow_219_fu_33033_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_221_fu_33211_p3 = ((overflow_220_fu_33182_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_222_fu_33360_p3 = ((overflow_221_fu_33331_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_223_fu_33509_p3 = ((overflow_222_fu_33480_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_224_fu_33534_p3 = ((overflow_223_reg_43330[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_225_fu_37176_p3 = ((overflow_224_fu_37147_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_226_fu_37300_p3 = ((overflow_225_fu_37271_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_227_fu_37425_p3 = ((overflow_226_fu_37396_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_228_fu_37550_p3 = ((overflow_227_fu_37521_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_229_fu_37675_p3 = ((overflow_228_fu_37646_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_230_fu_37800_p3 = ((overflow_229_fu_37771_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_231_fu_37925_p3 = ((overflow_230_fu_37896_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_232_fu_38050_p3 = ((overflow_231_fu_38021_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_233_fu_38175_p3 = ((overflow_232_fu_38146_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_234_fu_38320_p3 = ((overflow_233_fu_38291_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_235_fu_38469_p3 = ((overflow_234_fu_38440_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_236_fu_38618_p3 = ((overflow_235_fu_38589_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_237_fu_38767_p3 = ((overflow_236_fu_38738_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_238_fu_38916_p3 = ((overflow_237_fu_38887_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_239_fu_39065_p3 = ((overflow_238_fu_39036_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_240_fu_39214_p3 = ((overflow_239_fu_39185_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_241_fu_39239_p3 = ((overflow_240_reg_44007[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_242_fu_39380_p3 = ((overflow_241_fu_39351_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_fu_19069_p3 = ((overflow_fu_19040_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln350_100_fu_29466_p3 = ((underflow_262_fu_29434_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_685_fu_29403_p2);

assign select_ln350_101_fu_29564_p3 = ((underflow_263_fu_29532_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_687_fu_29502_p2);

assign select_ln350_102_fu_29664_p3 = ((underflow_264_fu_29632_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_689_fu_29601_p2);

assign select_ln350_103_fu_29764_p3 = ((underflow_265_fu_29732_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_691_fu_29701_p2);

assign select_ln350_104_fu_29864_p3 = ((underflow_266_fu_29832_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_693_fu_29801_p2);

assign select_ln350_105_fu_29964_p3 = ((underflow_267_fu_29932_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_695_fu_29901_p2);

assign select_ln350_106_fu_30064_p3 = ((underflow_268_fu_30032_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_697_fu_30001_p2);

assign select_ln350_107_fu_30166_p3 = ((underflow_269_fu_30134_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_699_fu_30102_p2);

assign select_ln350_108_fu_30268_p3 = ((underflow_270_fu_30236_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_701_fu_30204_p2);

assign select_ln350_109_fu_30370_p3 = ((underflow_271_fu_30338_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_703_fu_30306_p2);

assign select_ln350_110_fu_30472_p3 = ((underflow_272_fu_30440_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_705_fu_30408_p2);

assign select_ln350_111_fu_30574_p3 = ((underflow_273_fu_30542_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_707_fu_30510_p2);

assign select_ln350_112_fu_30676_p3 = ((underflow_274_fu_30644_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_709_fu_30612_p2);

assign select_ln350_113_fu_30778_p3 = ((underflow_275_fu_30746_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_711_fu_30714_p2);

assign select_ln350_114_fu_30880_p3 = ((underflow_276_fu_30848_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_713_fu_30816_p2);

assign select_ln350_115_fu_30982_p3 = ((underflow_277_fu_30950_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_715_fu_30918_p2);

assign select_ln350_116_fu_34761_p3 = ((underflow_278_fu_34733_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_717_reg_43347);

assign select_ln350_117_fu_34819_p3 = ((underflow_279_fu_34791_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_719_reg_43367);

assign select_ln350_118_fu_34877_p3 = ((underflow_280_fu_34849_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_721_reg_43387);

assign select_ln350_119_fu_34935_p3 = ((underflow_281_fu_34907_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_723_reg_43407);

assign select_ln350_120_fu_34993_p3 = ((underflow_282_fu_34965_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_725_reg_43427);

assign select_ln350_121_fu_35051_p3 = ((underflow_283_fu_35023_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_727_reg_43447);

assign select_ln350_122_fu_35109_p3 = ((underflow_284_fu_35081_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_729_reg_43467);

assign select_ln350_123_fu_35167_p3 = ((underflow_285_fu_35139_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_731_reg_43487);

assign select_ln350_124_fu_35225_p3 = ((underflow_286_fu_35197_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_733_reg_43507);

assign select_ln350_125_fu_35326_p3 = ((underflow_287_fu_35294_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_735_fu_35262_p2);

assign select_ln350_126_fu_35428_p3 = ((underflow_288_fu_35396_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_737_fu_35364_p2);

assign select_ln350_127_fu_35530_p3 = ((underflow_289_fu_35498_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_739_fu_35466_p2);

assign select_ln350_128_fu_35632_p3 = ((underflow_290_fu_35600_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_741_fu_35568_p2);

assign select_ln350_129_fu_35734_p3 = ((underflow_291_fu_35702_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_743_fu_35670_p2);

assign select_ln350_130_fu_35836_p3 = ((underflow_292_fu_35804_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_745_fu_35772_p2);

assign select_ln350_131_fu_35938_p3 = ((underflow_293_fu_35906_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_747_fu_35874_p2);

assign select_ln350_132_fu_36040_p3 = ((underflow_294_fu_36008_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_749_fu_35976_p2);

assign select_ln350_133_fu_36142_p3 = ((underflow_295_fu_36110_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_751_fu_36078_p2);

assign select_ln350_134_fu_36244_p3 = ((underflow_296_fu_36212_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_753_fu_36180_p2);

assign select_ln350_135_fu_36346_p3 = ((underflow_297_fu_36314_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_755_fu_36282_p2);

assign select_ln350_136_fu_36448_p3 = ((underflow_298_fu_36416_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_757_fu_36384_p2);

assign select_ln350_137_fu_36550_p3 = ((underflow_299_fu_36518_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_759_fu_36486_p2);

assign select_ln350_138_fu_36652_p3 = ((underflow_300_fu_36620_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_761_fu_36588_p2);

assign select_ln350_139_fu_36754_p3 = ((underflow_301_fu_36722_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_763_fu_36690_p2);

assign select_ln350_140_fu_36856_p3 = ((underflow_302_fu_36824_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_765_fu_36792_p2);

assign select_ln350_141_fu_36958_p3 = ((underflow_303_fu_36926_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_767_fu_36894_p2);

assign select_ln350_142_fu_37060_p3 = ((underflow_304_fu_37028_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_769_fu_36996_p2);

assign select_ln350_143_fu_39486_p3 = ((underflow_305_fu_39454_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_771_fu_39423_p2);

assign select_ln350_144_fu_39586_p3 = ((underflow_306_fu_39554_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_773_fu_39523_p2);

assign select_ln350_145_fu_39686_p3 = ((underflow_307_fu_39654_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_775_fu_39623_p2);

assign select_ln350_146_fu_39786_p3 = ((underflow_308_fu_39754_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_777_fu_39723_p2);

assign select_ln350_147_fu_39886_p3 = ((underflow_309_fu_39854_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_779_fu_39823_p2);

assign select_ln350_148_fu_39986_p3 = ((underflow_310_fu_39954_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_781_fu_39923_p2);

assign select_ln350_149_fu_40086_p3 = ((underflow_311_fu_40054_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_783_fu_40023_p2);

assign select_ln350_150_fu_40186_p3 = ((underflow_312_fu_40154_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_785_fu_40123_p2);

assign select_ln350_151_fu_40286_p3 = ((underflow_313_fu_40254_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_787_fu_40223_p2);

assign select_ln350_152_fu_40388_p3 = ((underflow_314_fu_40356_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_789_fu_40324_p2);

assign select_ln350_153_fu_40490_p3 = ((underflow_315_fu_40458_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_791_fu_40426_p2);

assign select_ln350_154_fu_40592_p3 = ((underflow_316_fu_40560_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_793_fu_40528_p2);

assign select_ln350_155_fu_40694_p3 = ((underflow_317_fu_40662_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_795_fu_40630_p2);

assign select_ln350_156_fu_40796_p3 = ((underflow_318_fu_40764_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_797_fu_40732_p2);

assign select_ln350_157_fu_40898_p3 = ((underflow_319_fu_40866_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_799_fu_40834_p2);

assign select_ln350_158_fu_41000_p3 = ((underflow_320_fu_40968_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_801_fu_40936_p2);

assign select_ln350_159_fu_41102_p3 = ((underflow_321_fu_41070_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_803_fu_41038_p2);

assign select_ln350_160_fu_41204_p3 = ((underflow_322_fu_41172_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_805_fu_41140_p2);

assign select_ln350_81_fu_23802_p3 = ((underflow_243_fu_23770_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_647_fu_23738_p2);

assign select_ln350_82_fu_23900_p3 = ((underflow_244_fu_23868_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_649_fu_23836_p2);

assign select_ln350_83_fu_23998_p3 = ((underflow_245_fu_23966_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_651_fu_23934_p2);

assign select_ln350_84_fu_24096_p3 = ((underflow_246_fu_24064_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_653_fu_24032_p2);

assign select_ln350_85_fu_24194_p3 = ((underflow_247_fu_24162_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_655_fu_24130_p2);

assign select_ln350_86_fu_24292_p3 = ((underflow_248_fu_24260_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_657_fu_24228_p2);

assign select_ln350_87_fu_24390_p3 = ((underflow_249_fu_24358_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_659_fu_24326_p2);

assign select_ln350_88_fu_24488_p3 = ((underflow_250_fu_24456_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_661_fu_24424_p2);

assign select_ln350_89_fu_24590_p3 = ((underflow_251_fu_24558_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_663_fu_24526_p2);

assign select_ln350_90_fu_24692_p3 = ((underflow_252_fu_24660_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_665_fu_24628_p2);

assign select_ln350_91_fu_24794_p3 = ((underflow_253_fu_24762_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_667_fu_24730_p2);

assign select_ln350_92_fu_24896_p3 = ((underflow_254_fu_24864_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_669_fu_24832_p2);

assign select_ln350_93_fu_24998_p3 = ((underflow_255_fu_24966_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_671_fu_24934_p2);

assign select_ln350_94_fu_25100_p3 = ((underflow_256_fu_25068_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_673_fu_25036_p2);

assign select_ln350_95_fu_25202_p3 = ((underflow_257_fu_25170_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_675_fu_25138_p2);

assign select_ln350_96_fu_25304_p3 = ((underflow_258_fu_25272_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_677_fu_25240_p2);

assign select_ln350_97_fu_25406_p3 = ((underflow_259_fu_25374_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_679_fu_25342_p2);

assign select_ln350_98_fu_29266_p3 = ((underflow_260_fu_29234_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_681_fu_29204_p2);

assign select_ln350_99_fu_29366_p3 = ((underflow_261_fu_29334_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_683_fu_29303_p2);

assign select_ln350_fu_23704_p3 = ((underflow_242_fu_23672_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_645_fu_23640_p2);

assign sext_ln1273_13_fu_18117_p1 = $signed(shl_ln1273_s_fu_18109_p3);

assign sext_ln1273_14_fu_22897_p1 = $signed(shl_ln1273_12_fu_22890_p3);

assign sext_ln1273_15_fu_22908_p1 = $signed(shl_ln1273_13_fu_22901_p3);

assign sext_ln1273_16_fu_27925_p1 = $signed(shl_ln1273_14_fu_27918_p3);

assign sext_ln1273_17_fu_27936_p1 = $signed(shl_ln1273_15_fu_27929_p3);

assign sext_ln1273_18_fu_28992_p1 = $signed(shl_ln1273_16_fu_28985_p3);

assign sext_ln1273_19_fu_29003_p1 = $signed(shl_ln1273_17_fu_28996_p3);

assign sext_ln1273_20_fu_34469_p1 = $signed(shl_ln1273_18_fu_34462_p3);

assign sext_ln1273_21_fu_34486_p1 = $signed(shl_ln1273_19_fu_34479_p3);

assign sext_ln1273_fu_18099_p1 = $signed(shl_ln_fu_18091_p3);

assign sext_ln70_46_fu_17254_p0 = p_read_int_reg;

assign sext_ln70_46_fu_17254_p1 = sext_ln70_46_fu_17254_p0;

assign sext_ln70_47_fu_17260_p0 = p_read_int_reg;

assign sext_ln70_47_fu_17260_p1 = sext_ln70_47_fu_17260_p0;

assign sext_ln70_48_fu_17266_p0 = p_read_int_reg;

assign sext_ln70_48_fu_17266_p1 = sext_ln70_48_fu_17266_p0;

assign sext_ln70_53_fu_17869_p0 = p_read1_int_reg;

assign sext_ln70_53_fu_17869_p1 = sext_ln70_53_fu_17869_p0;

assign sext_ln70_60_fu_18458_p0 = p_read2_int_reg;

assign sext_ln70_60_fu_18458_p1 = sext_ln70_60_fu_18458_p0;

assign sext_ln70_63_fu_22489_p1 = p_read_32_reg_41324;

assign sext_ln70_64_fu_22494_p1 = p_read_32_reg_41324;

assign sext_ln70_65_fu_22500_p1 = p_read_32_reg_41324;

assign sext_ln70_66_fu_23217_p1 = p_read_31_reg_41314;

assign sext_ln70_69_fu_23230_p1 = p_read_31_reg_41314;

assign sext_ln70_74_fu_27903_p1 = p_read_30_reg_41303_pp0_iter1_reg;

assign sext_ln70_75_fu_27908_p1 = p_read_30_reg_41303_pp0_iter1_reg;

assign sext_ln70_79_fu_28637_p1 = p_read_29_reg_41293_pp0_iter1_reg;

assign sext_ln70_80_fu_28644_p1 = p_read_29_reg_41293_pp0_iter1_reg;

assign sext_ln70_81_fu_33548_p1 = p_read_28_reg_41284_pp0_iter2_reg;

assign sext_ln70_84_fu_33561_p1 = p_read_28_reg_41284_pp0_iter2_reg;

assign sext_ln70_86_fu_34148_p1 = p_read_27_reg_41274_pp0_iter2_reg;

assign sext_ln70_87_fu_34154_p1 = p_read_27_reg_41274_pp0_iter2_reg;

assign sext_ln70_88_fu_34159_p1 = p_read_27_reg_41274_pp0_iter2_reg;

assign sext_ln813_153_fu_23720_p1 = rhs_81_fu_19208_p3;

assign sext_ln813_154_fu_23818_p1 = rhs_82_fu_19333_p3;

assign sext_ln813_155_fu_23916_p1 = rhs_83_fu_19458_p3;

assign sext_ln813_156_fu_24014_p1 = rhs_84_fu_19583_p3;

assign sext_ln813_157_fu_24112_p1 = rhs_85_fu_19708_p3;

assign sext_ln813_158_fu_24210_p1 = rhs_86_fu_19833_p3;

assign sext_ln813_159_fu_24308_p1 = rhs_87_fu_19958_p3;

assign sext_ln813_160_fu_24406_p1 = rhs_88_fu_20083_p3;

assign sext_ln813_161_fu_24504_p1 = lhs_fu_23712_p3;

assign sext_ln813_162_fu_24508_p1 = rhs_89_fu_20232_p3;

assign sext_ln813_163_fu_24606_p1 = lhs_72_fu_23810_p3;

assign sext_ln813_164_fu_24610_p1 = rhs_90_fu_20381_p3;

assign sext_ln813_165_fu_24708_p1 = lhs_73_fu_23908_p3;

assign sext_ln813_166_fu_24712_p1 = rhs_91_fu_20530_p3;

assign sext_ln813_167_fu_24810_p1 = lhs_74_fu_24006_p3;

assign sext_ln813_168_fu_24814_p1 = rhs_92_fu_20679_p3;

assign sext_ln813_169_fu_24912_p1 = lhs_75_fu_24104_p3;

assign sext_ln813_170_fu_24916_p1 = rhs_93_fu_20828_p3;

assign sext_ln813_171_fu_25014_p1 = lhs_76_fu_24202_p3;

assign sext_ln813_172_fu_25018_p1 = rhs_94_fu_20846_p3;

assign sext_ln813_173_fu_25116_p1 = lhs_77_fu_24300_p3;

assign sext_ln813_174_fu_25120_p1 = rhs_95_fu_20994_p3;

assign sext_ln813_175_fu_25218_p1 = lhs_78_fu_24398_p3;

assign sext_ln813_176_fu_25222_p1 = rhs_96_fu_21143_p3;

assign sext_ln813_177_fu_25320_p1 = lhs_79_fu_24496_p3;

assign sext_ln813_178_fu_25324_p1 = rhs_97_fu_21292_p3;

assign sext_ln813_179_fu_29184_p1 = lhs_80_reg_42776;

assign sext_ln813_180_fu_29187_p1 = rhs_98_reg_42135;

assign sext_ln813_181_fu_29282_p1 = lhs_81_reg_42782;

assign sext_ln813_182_fu_29285_p1 = rhs_99_fu_25432_p3;

assign sext_ln813_183_fu_29382_p1 = lhs_82_reg_42788;

assign sext_ln813_184_fu_29385_p1 = rhs_100_fu_25449_p3;

assign sext_ln813_185_fu_29482_p1 = lhs_83_reg_42794;

assign sext_ln813_186_fu_29485_p1 = rhs_101_reg_42171;

assign sext_ln813_187_fu_29580_p1 = lhs_84_reg_42800;

assign sext_ln813_188_fu_29583_p1 = rhs_102_fu_25466_p3;

assign sext_ln813_189_fu_29680_p1 = lhs_85_reg_42806;

assign sext_ln813_190_fu_29683_p1 = rhs_103_fu_25483_p3;

assign sext_ln813_191_fu_29780_p1 = lhs_86_reg_42812;

assign sext_ln813_192_fu_29783_p1 = rhs_104_fu_25500_p3;

assign sext_ln813_193_fu_29880_p1 = lhs_87_reg_42818;

assign sext_ln813_194_fu_29883_p1 = rhs_105_fu_25517_p3;

assign sext_ln813_195_fu_29980_p1 = lhs_88_reg_42824;

assign sext_ln813_196_fu_29983_p1 = rhs_106_fu_25534_p3;

assign sext_ln813_197_fu_30080_p1 = lhs_89_fu_29274_p3;

assign sext_ln813_198_fu_30084_p1 = rhs_107_fu_25658_p3;

assign sext_ln813_199_fu_30182_p1 = lhs_90_fu_29374_p3;

assign sext_ln813_200_fu_30186_p1 = rhs_108_fu_25783_p3;

assign sext_ln813_201_fu_30284_p1 = lhs_91_fu_29474_p3;

assign sext_ln813_202_fu_30288_p1 = rhs_109_fu_25908_p3;

assign sext_ln813_203_fu_30386_p1 = lhs_92_fu_29572_p3;

assign sext_ln813_204_fu_30390_p1 = rhs_110_fu_26033_p3;

assign sext_ln813_205_fu_30488_p1 = lhs_93_fu_29672_p3;

assign sext_ln813_206_fu_30492_p1 = rhs_111_fu_26158_p3;

assign sext_ln813_207_fu_30590_p1 = lhs_94_fu_29772_p3;

assign sext_ln813_208_fu_30594_p1 = rhs_112_fu_26283_p3;

assign sext_ln813_209_fu_30692_p1 = lhs_95_fu_29872_p3;

assign sext_ln813_210_fu_30696_p1 = rhs_113_fu_26301_p3;

assign sext_ln813_211_fu_30794_p1 = lhs_96_fu_29972_p3;

assign sext_ln813_212_fu_30798_p1 = rhs_114_fu_26425_p3;

assign sext_ln813_213_fu_30896_p1 = lhs_97_fu_30072_p3;

assign sext_ln813_214_fu_30900_p1 = rhs_115_fu_26550_p3;

assign sext_ln813_215_fu_30998_p1 = lhs_98_fu_30174_p3;

assign sext_ln813_216_fu_31002_p1 = rhs_116_fu_26695_p3;

assign sext_ln813_217_fu_31034_p1 = lhs_99_fu_30276_p3;

assign sext_ln813_218_fu_31038_p1 = rhs_117_fu_26844_p3;

assign sext_ln813_219_fu_31070_p1 = lhs_100_fu_30378_p3;

assign sext_ln813_220_fu_31074_p1 = rhs_118_fu_26993_p3;

assign sext_ln813_221_fu_31106_p1 = lhs_101_fu_30480_p3;

assign sext_ln813_222_fu_31110_p1 = rhs_119_fu_27142_p3;

assign sext_ln813_223_fu_31142_p1 = lhs_102_fu_30582_p3;

assign sext_ln813_224_fu_31146_p1 = rhs_120_fu_27291_p3;

assign sext_ln813_225_fu_31178_p1 = lhs_103_fu_30684_p3;

assign sext_ln813_226_fu_31182_p1 = rhs_121_fu_27440_p3;

assign sext_ln813_227_fu_31214_p1 = lhs_104_fu_30786_p3;

assign sext_ln813_228_fu_31218_p1 = rhs_122_fu_27589_p3;

assign sext_ln813_229_fu_31250_p1 = lhs_105_fu_30888_p3;

assign sext_ln813_230_fu_31254_p1 = rhs_123_fu_27738_p3;

assign sext_ln813_231_fu_31286_p1 = lhs_106_fu_30990_p3;

assign sext_ln813_232_fu_31290_p1 = rhs_124_fu_27887_p3;

assign sext_ln813_233_fu_35240_p1 = lhs_107_fu_34768_p3;

assign sext_ln813_234_fu_35244_p1 = rhs_125_fu_31332_p3;

assign sext_ln813_235_fu_35342_p1 = lhs_108_fu_34826_p3;

assign sext_ln813_236_fu_35346_p1 = rhs_126_fu_31456_p3;

assign sext_ln813_237_fu_35444_p1 = lhs_109_fu_34884_p3;

assign sext_ln813_238_fu_35448_p1 = rhs_127_fu_31581_p3;

assign sext_ln813_239_fu_35546_p1 = lhs_110_fu_34942_p3;

assign sext_ln813_240_fu_35550_p1 = rhs_128_fu_31706_p3;

assign sext_ln813_241_fu_35648_p1 = lhs_111_fu_35000_p3;

assign sext_ln813_242_fu_35652_p1 = rhs_129_fu_31831_p3;

assign sext_ln813_243_fu_35750_p1 = lhs_112_fu_35058_p3;

assign sext_ln813_244_fu_35754_p1 = rhs_130_fu_31956_p3;

assign sext_ln813_245_fu_35852_p1 = lhs_113_fu_35116_p3;

assign sext_ln813_246_fu_35856_p1 = rhs_131_fu_32081_p3;

assign sext_ln813_247_fu_35954_p1 = lhs_114_fu_35174_p3;

assign sext_ln813_248_fu_35958_p1 = rhs_132_fu_32206_p3;

assign sext_ln813_249_fu_36056_p1 = lhs_115_fu_35232_p3;

assign sext_ln813_250_fu_36060_p1 = rhs_133_fu_32331_p3;

assign sext_ln813_251_fu_36158_p1 = lhs_116_fu_35334_p3;

assign sext_ln813_252_fu_36162_p1 = rhs_134_fu_32480_p3;

assign sext_ln813_253_fu_36260_p1 = lhs_117_fu_35436_p3;

assign sext_ln813_254_fu_36264_p1 = rhs_135_fu_32629_p3;

assign sext_ln813_255_fu_36362_p1 = lhs_118_fu_35538_p3;

assign sext_ln813_256_fu_36366_p1 = rhs_136_fu_32778_p3;

assign sext_ln813_257_fu_36464_p1 = lhs_119_fu_35640_p3;

assign sext_ln813_258_fu_36468_p1 = rhs_137_fu_32927_p3;

assign sext_ln813_259_fu_36566_p1 = lhs_120_fu_35742_p3;

assign sext_ln813_260_fu_36570_p1 = rhs_138_fu_33076_p3;

assign sext_ln813_261_fu_36668_p1 = lhs_121_fu_35844_p3;

assign sext_ln813_262_fu_36672_p1 = rhs_139_fu_33225_p3;

assign sext_ln813_263_fu_36770_p1 = lhs_122_fu_35946_p3;

assign sext_ln813_264_fu_36774_p1 = rhs_140_fu_33374_p3;

assign sext_ln813_265_fu_36872_p1 = lhs_123_fu_36048_p3;

assign sext_ln813_266_fu_36876_p1 = rhs_141_fu_33523_p3;

assign sext_ln813_267_fu_36974_p1 = lhs_124_fu_36150_p3;

assign sext_ln813_268_fu_36978_p1 = rhs_142_fu_33541_p3;

assign sext_ln813_269_fu_39402_p1 = lhs_125_reg_44046;

assign sext_ln813_270_fu_39405_p1 = rhs_143_fu_37190_p3;

assign sext_ln813_271_fu_39502_p1 = lhs_126_reg_44052;

assign sext_ln813_272_fu_39505_p1 = rhs_144_fu_37314_p3;

assign sext_ln813_273_fu_39602_p1 = lhs_127_reg_44058;

assign sext_ln813_274_fu_39605_p1 = rhs_145_fu_37439_p3;

assign sext_ln813_275_fu_39702_p1 = lhs_128_reg_44064;

assign sext_ln813_276_fu_39705_p1 = rhs_146_fu_37564_p3;

assign sext_ln813_277_fu_39802_p1 = lhs_129_reg_44070;

assign sext_ln813_278_fu_39805_p1 = rhs_147_fu_37689_p3;

assign sext_ln813_279_fu_39902_p1 = lhs_130_reg_44076;

assign sext_ln813_280_fu_39905_p1 = rhs_148_fu_37814_p3;

assign sext_ln813_281_fu_40002_p1 = lhs_131_reg_44082;

assign sext_ln813_282_fu_40005_p1 = rhs_149_fu_37939_p3;

assign sext_ln813_283_fu_40102_p1 = lhs_132_reg_44088;

assign sext_ln813_284_fu_40105_p1 = rhs_150_fu_38064_p3;

assign sext_ln813_285_fu_40202_p1 = lhs_133_reg_44094;

assign sext_ln813_286_fu_40205_p1 = rhs_151_fu_38189_p3;

assign sext_ln813_287_fu_40302_p1 = lhs_134_fu_39494_p3;

assign sext_ln813_288_fu_40306_p1 = rhs_152_fu_38334_p3;

assign sext_ln813_289_fu_40404_p1 = lhs_135_fu_39594_p3;

assign sext_ln813_290_fu_40408_p1 = rhs_153_fu_38483_p3;

assign sext_ln813_291_fu_40506_p1 = lhs_136_fu_39694_p3;

assign sext_ln813_292_fu_40510_p1 = rhs_154_fu_38632_p3;

assign sext_ln813_293_fu_40608_p1 = lhs_137_fu_39794_p3;

assign sext_ln813_294_fu_40612_p1 = rhs_155_fu_38781_p3;

assign sext_ln813_295_fu_40710_p1 = lhs_138_fu_39894_p3;

assign sext_ln813_296_fu_40714_p1 = rhs_156_fu_38930_p3;

assign sext_ln813_297_fu_40812_p1 = lhs_139_fu_39994_p3;

assign sext_ln813_298_fu_40816_p1 = rhs_157_fu_39079_p3;

assign sext_ln813_299_fu_40914_p1 = lhs_140_fu_40094_p3;

assign sext_ln813_300_fu_40918_p1 = rhs_158_fu_39228_p3;

assign sext_ln813_301_fu_41016_p1 = lhs_141_fu_40194_p3;

assign sext_ln813_302_fu_41020_p1 = rhs_159_fu_39246_p3;

assign sext_ln813_303_fu_41118_p1 = lhs_142_fu_40294_p3;

assign sext_ln813_304_fu_41122_p1 = rhs_160_fu_39394_p3;

assign sext_ln813_fu_23622_p1 = rhs_fu_19083_p3;

assign sext_ln818_1_fu_26558_p1 = $signed(p_Val2_510_reg_42521);

assign sext_ln818_2_fu_33590_p1 = $signed(p_Val2_591_fu_33580_p4);

assign sext_ln818_3_fu_38197_p1 = $signed(p_Val2_618_reg_43805);

assign sext_ln818_fu_21300_p1 = $signed(p_Val2_456_reg_41865);

assign sext_ln823_100_fu_22231_p1 = $signed(p_Val2_477_reg_42068);

assign sext_ln823_101_fu_22360_p1 = $signed(p_Val2_480_reg_42097);

assign sext_ln823_102_fu_22524_p1 = $signed(p_Val2_483_fu_22514_p4);

assign sext_ln823_103_fu_22588_p1 = $signed(p_Val2_486_fu_22578_p4);

assign sext_ln823_104_fu_22652_p1 = $signed(p_Val2_489_fu_22642_p4);

assign sext_ln823_105_fu_22716_p1 = $signed(p_Val2_492_fu_22706_p4);

assign sext_ln823_106_fu_22780_p1 = $signed(p_Val2_495_fu_22770_p4);

assign sext_ln823_107_fu_22844_p1 = $signed(p_Val2_498_fu_22834_p4);

assign sext_ln823_108_fu_22936_p1 = $signed(p_Val2_501_fu_22926_p4);

assign sext_ln823_109_fu_23107_p1 = $signed(p_Val2_504_fu_23097_p4);

assign sext_ln823_110_fu_23171_p1 = $signed(p_Val2_507_fu_23161_p4);

assign sext_ln823_111_fu_26703_p1 = $signed(p_Val2_513_reg_42550);

assign sext_ln823_112_fu_26852_p1 = $signed(p_Val2_516_reg_42579);

assign sext_ln823_113_fu_27001_p1 = $signed(p_Val2_519_reg_42608);

assign sext_ln823_114_fu_27150_p1 = $signed(p_Val2_522_reg_42637);

assign sext_ln823_115_fu_27299_p1 = $signed(p_Val2_525_reg_42666);

assign sext_ln823_116_fu_27448_p1 = $signed(p_Val2_528_reg_42695);

assign sext_ln823_117_fu_27597_p1 = $signed(p_Val2_531_reg_42724);

assign sext_ln823_118_fu_27746_p1 = $signed(p_Val2_534_reg_42753);

assign sext_ln823_119_fu_27964_p1 = $signed(p_Val2_537_fu_27954_p4);

assign sext_ln823_120_fu_28135_p1 = $signed(p_Val2_540_fu_28125_p4);

assign sext_ln823_121_fu_28199_p1 = $signed(p_Val2_543_fu_28189_p4);

assign sext_ln823_122_fu_28263_p1 = $signed(p_Val2_546_fu_28253_p4);

assign sext_ln823_123_fu_28327_p1 = $signed(p_Val2_549_fu_28317_p4);

assign sext_ln823_124_fu_28391_p1 = $signed(p_Val2_552_fu_28381_p4);

assign sext_ln823_125_fu_28455_p1 = $signed(p_Val2_555_fu_28445_p4);

assign sext_ln823_126_fu_28519_p1 = $signed(p_Val2_558_fu_28509_p4);

assign sext_ln823_127_fu_28583_p1 = $signed(p_Val2_561_fu_28573_p4);

assign sext_ln823_128_fu_32339_p1 = $signed(p_Val2_564_reg_43099);

assign sext_ln823_129_fu_32488_p1 = $signed(p_Val2_567_reg_43128);

assign sext_ln823_130_fu_32637_p1 = $signed(p_Val2_570_reg_43157);

assign sext_ln823_131_fu_32786_p1 = $signed(p_Val2_573_reg_43186);

assign sext_ln823_132_fu_32935_p1 = $signed(p_Val2_576_reg_43215);

assign sext_ln823_133_fu_33084_p1 = $signed(p_Val2_579_reg_43244);

assign sext_ln823_134_fu_33233_p1 = $signed(p_Val2_582_reg_43273);

assign sext_ln823_135_fu_33382_p1 = $signed(p_Val2_585_reg_43302);

assign sext_ln823_136_fu_29031_p1 = $signed(p_Val2_588_fu_29021_p4);

assign sext_ln823_137_fu_33654_p1 = $signed(p_Val2_594_fu_33644_p4);

assign sext_ln823_138_fu_33718_p1 = $signed(p_Val2_597_fu_33708_p4);

assign sext_ln823_139_fu_33782_p1 = $signed(p_Val2_600_fu_33772_p4);

assign sext_ln823_140_fu_33846_p1 = $signed(p_Val2_603_fu_33836_p4);

assign sext_ln823_141_fu_33910_p1 = $signed(p_Val2_606_fu_33900_p4);

assign sext_ln823_142_fu_33974_p1 = $signed(p_Val2_609_fu_33964_p4);

assign sext_ln823_143_fu_34038_p1 = $signed(p_Val2_612_fu_34028_p4);

assign sext_ln823_144_fu_34102_p1 = $signed(p_Val2_615_fu_34092_p4);

assign sext_ln823_145_fu_38342_p1 = $signed(p_Val2_621_reg_43834);

assign sext_ln823_146_fu_38491_p1 = $signed(p_Val2_624_reg_43863);

assign sext_ln823_147_fu_38640_p1 = $signed(p_Val2_627_reg_43892);

assign sext_ln823_148_fu_38789_p1 = $signed(p_Val2_630_reg_43921);

assign sext_ln823_149_fu_38938_p1 = $signed(p_Val2_633_reg_43950);

assign sext_ln823_150_fu_39087_p1 = $signed(p_Val2_636_reg_43979);

assign sext_ln823_151_fu_34514_p1 = $signed(p_Val2_639_fu_34504_p4);

assign sext_ln823_152_fu_39253_p1 = $signed(p_Val2_642_reg_44023);

assign sext_ln823_78_fu_17355_p1 = $signed(p_Val2_405_fu_17345_p4);

assign sext_ln823_79_fu_17419_p1 = $signed(p_Val2_408_fu_17409_p4);

assign sext_ln823_80_fu_17483_p1 = $signed(p_Val2_411_fu_17473_p4);

assign sext_ln823_81_fu_17547_p1 = $signed(p_Val2_414_fu_17537_p4);

assign sext_ln823_82_fu_17611_p1 = $signed(p_Val2_417_fu_17601_p4);

assign sext_ln823_83_fu_17675_p1 = $signed(p_Val2_420_fu_17665_p4);

assign sext_ln823_84_fu_17739_p1 = $signed(p_Val2_423_fu_17729_p4);

assign sext_ln823_85_fu_17803_p1 = $signed(p_Val2_426_fu_17793_p4);

assign sext_ln823_86_fu_20091_p1 = $signed(p_Val2_429_reg_41618);

assign sext_ln823_87_fu_20240_p1 = $signed(p_Val2_432_reg_41647);

assign sext_ln823_88_fu_20389_p1 = $signed(p_Val2_435_reg_41676);

assign sext_ln823_89_fu_20538_p1 = $signed(p_Val2_438_reg_41705);

assign sext_ln823_90_fu_20687_p1 = $signed(p_Val2_441_reg_41734);

assign sext_ln823_91_fu_18145_p1 = $signed(p_Val2_444_fu_18135_p4);

assign sext_ln823_92_fu_20853_p1 = $signed(p_Val2_447_reg_41778);

assign sext_ln823_93_fu_21002_p1 = $signed(p_Val2_450_reg_41807);

assign sext_ln823_94_fu_21151_p1 = $signed(p_Val2_453_reg_41836);

assign sext_ln823_95_fu_21445_p1 = $signed(p_Val2_459_reg_41894);

assign sext_ln823_96_fu_21574_p1 = $signed(p_Val2_462_reg_41923);

assign sext_ln823_97_fu_21844_p1 = $signed(p_Val2_468_reg_41981);

assign sext_ln823_98_fu_21973_p1 = $signed(p_Val2_471_reg_42010);

assign sext_ln823_99_fu_22102_p1 = $signed(p_Val2_474_reg_42039);

assign sext_ln823_fu_17291_p1 = $signed(p_Val2_402_fu_17281_p4);

assign sext_ln856_100_fu_25507_p1 = p_Val2_478_reg_42222;

assign sext_ln856_101_fu_25524_p1 = p_Val2_481_reg_42237;

assign sext_ln856_102_fu_25541_p1 = p_Val2_484_reg_42264;

assign sext_ln856_103_fu_25666_p1 = p_Val2_487_reg_42295;

assign sext_ln856_104_fu_25791_p1 = p_Val2_490_reg_42326;

assign sext_ln856_105_fu_25916_p1 = p_Val2_493_reg_42357;

assign sext_ln856_106_fu_26041_p1 = p_Val2_496_reg_42388;

assign sext_ln856_107_fu_26166_p1 = p_Val2_499_reg_42419;

assign sext_ln856_108_fu_26291_p1 = p_Val2_502_reg_42438;

assign sext_ln856_109_fu_26308_p1 = p_Val2_505_reg_42465;

assign sext_ln856_110_fu_26433_p1 = p_Val2_508_reg_42496;

assign sext_ln856_111_fu_26715_p1 = p_Val2_514_fu_26709_p2;

assign sext_ln856_112_fu_26864_p1 = p_Val2_517_fu_26858_p2;

assign sext_ln856_113_fu_27013_p1 = p_Val2_520_fu_27007_p2;

assign sext_ln856_114_fu_27162_p1 = p_Val2_523_fu_27156_p2;

assign sext_ln856_115_fu_27311_p1 = p_Val2_526_fu_27305_p2;

assign sext_ln856_116_fu_27460_p1 = p_Val2_529_fu_27454_p2;

assign sext_ln856_117_fu_27609_p1 = p_Val2_532_fu_27603_p2;

assign sext_ln856_118_fu_27758_p1 = p_Val2_535_fu_27752_p2;

assign sext_ln856_119_fu_31322_p1 = p_Val2_538_reg_42830;

assign sext_ln856_120_fu_31339_p1 = p_Val2_541_reg_42857;

assign sext_ln856_121_fu_31464_p1 = p_Val2_544_reg_42888;

assign sext_ln856_122_fu_31589_p1 = p_Val2_547_reg_42919;

assign sext_ln856_123_fu_31714_p1 = p_Val2_550_reg_42950;

assign sext_ln856_124_fu_31839_p1 = p_Val2_553_reg_42981;

assign sext_ln856_125_fu_31964_p1 = p_Val2_556_reg_43012;

assign sext_ln856_126_fu_32089_p1 = p_Val2_559_reg_43043;

assign sext_ln856_127_fu_32214_p1 = p_Val2_562_reg_43074;

assign sext_ln856_128_fu_32351_p1 = p_Val2_565_fu_32345_p2;

assign sext_ln856_129_fu_32500_p1 = p_Val2_568_fu_32494_p2;

assign sext_ln856_130_fu_32649_p1 = p_Val2_571_fu_32643_p2;

assign sext_ln856_131_fu_32798_p1 = p_Val2_574_fu_32792_p2;

assign sext_ln856_132_fu_32947_p1 = p_Val2_577_fu_32941_p2;

assign sext_ln856_133_fu_33096_p1 = p_Val2_580_fu_33090_p2;

assign sext_ln856_134_fu_33245_p1 = p_Val2_583_fu_33239_p2;

assign sext_ln856_135_fu_33394_p1 = p_Val2_586_fu_33388_p2;

assign sext_ln856_136_fu_33531_p1 = p_Val2_589_reg_43325;

assign sext_ln856_137_fu_37197_p1 = p_Val2_595_reg_43563;

assign sext_ln856_138_fu_37322_p1 = p_Val2_598_reg_43594;

assign sext_ln856_139_fu_37447_p1 = p_Val2_601_reg_43625;

assign sext_ln856_140_fu_37572_p1 = p_Val2_604_reg_43656;

assign sext_ln856_141_fu_37697_p1 = p_Val2_607_reg_43687;

assign sext_ln856_142_fu_37822_p1 = p_Val2_610_reg_43718;

assign sext_ln856_143_fu_37947_p1 = p_Val2_613_reg_43749;

assign sext_ln856_144_fu_38072_p1 = p_Val2_616_reg_43780;

assign sext_ln856_145_fu_38354_p1 = p_Val2_622_fu_38348_p2;

assign sext_ln856_146_fu_38503_p1 = p_Val2_625_fu_38497_p2;

assign sext_ln856_147_fu_38652_p1 = p_Val2_628_fu_38646_p2;

assign sext_ln856_148_fu_38801_p1 = p_Val2_631_fu_38795_p2;

assign sext_ln856_149_fu_38950_p1 = p_Val2_634_fu_38944_p2;

assign sext_ln856_150_fu_39099_p1 = p_Val2_637_fu_39093_p2;

assign sext_ln856_151_fu_39236_p1 = p_Val2_640_reg_44002;

assign sext_ln856_152_fu_39265_p1 = p_Val2_643_fu_39259_p2;

assign sext_ln856_78_fu_19091_p1 = p_Val2_406_reg_41376;

assign sext_ln856_79_fu_19216_p1 = p_Val2_409_reg_41407;

assign sext_ln856_80_fu_19341_p1 = p_Val2_412_reg_41438;

assign sext_ln856_81_fu_19466_p1 = p_Val2_415_reg_41469;

assign sext_ln856_82_fu_19591_p1 = p_Val2_418_reg_41500;

assign sext_ln856_83_fu_19716_p1 = p_Val2_421_reg_41531;

assign sext_ln856_84_fu_19841_p1 = p_Val2_424_reg_41562;

assign sext_ln856_85_fu_19966_p1 = p_Val2_427_reg_41593;

assign sext_ln856_86_fu_20103_p1 = p_Val2_430_fu_20097_p2;

assign sext_ln856_87_fu_20252_p1 = p_Val2_433_fu_20246_p2;

assign sext_ln856_88_fu_20401_p1 = p_Val2_436_fu_20395_p2;

assign sext_ln856_89_fu_20550_p1 = p_Val2_439_fu_20544_p2;

assign sext_ln856_90_fu_20699_p1 = p_Val2_442_fu_20693_p2;

assign sext_ln856_91_fu_20836_p1 = p_Val2_445_reg_41757;

assign sext_ln856_92_fu_20865_p1 = p_Val2_448_fu_20859_p2;

assign sext_ln856_93_fu_21014_p1 = p_Val2_451_fu_21008_p2;

assign sext_ln856_94_fu_21163_p1 = p_Val2_454_fu_21157_p2;

assign sext_ln856_95_fu_25422_p1 = p_Val2_460_reg_42141;

assign sext_ln856_96_fu_25439_p1 = p_Val2_463_reg_42156;

assign sext_ln856_97_fu_25456_p1 = p_Val2_469_reg_42177;

assign sext_ln856_98_fu_25473_p1 = p_Val2_472_reg_42192;

assign sext_ln856_99_fu_25490_p1 = p_Val2_475_reg_42207;

assign sext_ln856_fu_18966_p1 = p_Val2_403_reg_41345;

assign shl_ln1273_12_fu_22890_p3 = {{p_read_32_reg_41324}, {6'd0}};

assign shl_ln1273_13_fu_22901_p3 = {{p_read_32_reg_41324}, {1'd0}};

assign shl_ln1273_14_fu_27918_p3 = {{p_read_30_reg_41303_pp0_iter1_reg}, {8'd0}};

assign shl_ln1273_15_fu_27929_p3 = {{p_read_30_reg_41303_pp0_iter1_reg}, {1'd0}};

assign shl_ln1273_16_fu_28985_p3 = {{p_read_29_reg_41293_pp0_iter1_reg}, {8'd0}};

assign shl_ln1273_17_fu_28996_p3 = {{p_read_29_reg_41293_pp0_iter1_reg}, {5'd0}};

assign shl_ln1273_18_fu_34462_p3 = {{p_read_27_reg_41274_pp0_iter2_reg}, {3'd0}};

assign shl_ln1273_19_fu_34479_p3 = {{p_read_27_reg_41274_pp0_iter2_reg}, {1'd0}};

assign shl_ln1273_s_fu_18109_p1 = p_read1_int_reg;

assign shl_ln1273_s_fu_18109_p3 = {{shl_ln1273_s_fu_18109_p1}, {1'd0}};

assign shl_ln_fu_18091_p1 = p_read1_int_reg;

assign shl_ln_fu_18091_p3 = {{shl_ln_fu_18091_p1}, {7'd0}};

assign sub_ln1273_10_fu_34473_p2 = ($signed(36'd0) - $signed(sext_ln1273_20_fu_34469_p1));

assign sub_ln1273_fu_18103_p2 = ($signed(40'd0) - $signed(sext_ln1273_fu_18099_p1));

assign sub_ln823_2_fu_18914_p2 = (trunc_ln1273_4_fu_18906_p3 - trunc_ln1273_3_fu_18894_p3);

assign sub_ln823_3_fu_18952_p2 = (trunc_ln1273_6_fu_18944_p3 - trunc_ln1273_5_fu_18932_p3);

assign sub_ln823_fu_18876_p2 = (trunc_ln1273_2_fu_18868_p3 - trunc_ln5_fu_18856_p3);

assign tmp_1002_fu_33284_p3 = r_V_137_reg_15603[32'd40];

assign tmp_1008_fu_33433_p3 = r_V_138_reg_15607[32'd41];

assign tmp_1014_fu_29098_p3 = r_V_139_fu_29007_p2[32'd40];

assign tmp_1017_fu_33602_p3 = r_V_140_fu_481_p2[32'd23];

assign tmp_1020_fu_37101_p3 = r_V_140_reg_17175[32'd54];

assign tmp_1023_fu_33666_p3 = r_V_141_fu_541_p2[32'd23];

assign tmp_1026_fu_37225_p3 = r_V_141_reg_17179[32'd43];

assign tmp_1029_fu_33730_p3 = r_V_142_fu_492_p2[32'd23];

assign tmp_1032_fu_37350_p3 = r_V_142_reg_17183[32'd42];

assign tmp_1035_fu_33794_p3 = r_V_143_fu_540_p2[32'd23];

assign tmp_1038_fu_37475_p3 = r_V_143_reg_17187[32'd49];

assign tmp_1041_fu_33858_p3 = r_V_144_fu_490_p2[32'd23];

assign tmp_1044_fu_37600_p3 = r_V_144_reg_17191[32'd48];

assign tmp_1047_fu_33922_p3 = r_V_145_fu_476_p2[32'd23];

assign tmp_1050_fu_37725_p3 = r_V_145_reg_17195[32'd43];

assign tmp_1053_fu_33986_p3 = r_V_146_fu_514_p2[32'd23];

assign tmp_1056_fu_37850_p3 = r_V_146_reg_17199[32'd43];

assign tmp_1059_fu_34050_p3 = r_V_147_fu_508_p2[32'd23];

assign tmp_1062_fu_37975_p3 = r_V_147_reg_17203[32'd43];

assign tmp_1065_fu_34114_p3 = r_V_148_fu_518_p2[32'd23];

assign tmp_1068_fu_38100_p3 = r_V_148_reg_17207[32'd48];

assign tmp_1074_fu_38244_p3 = r_V_149_reg_17211[32'd54];

assign tmp_1080_fu_38393_p3 = r_V_150_reg_17215[32'd41];

assign tmp_1086_fu_38542_p3 = r_V_151_reg_17219[32'd43];

assign tmp_1092_fu_38691_p3 = r_V_152_reg_17223[32'd49];

assign tmp_1098_fu_38840_p3 = r_V_153_reg_17227[32'd49];

assign tmp_1104_fu_38989_p3 = r_V_154_reg_17231[32'd41];

assign tmp_1110_fu_39138_p3 = r_V_155_reg_17235[32'd43];

assign tmp_1113_fu_34526_p3 = r_V_156_fu_34490_p2[32'd23];

assign tmp_1116_fu_34590_p3 = r_V_156_fu_34490_p2[32'd35];

assign tmp_1122_fu_39304_p3 = r_V_157_reg_17239[32'd49];

assign tmp_642_fu_18994_p3 = r_V_reg_9071[32'd41];

assign tmp_645_fu_17367_p3 = r_V_78_fu_527_p2[32'd23];

assign tmp_648_fu_19119_p3 = r_V_78_reg_9075[32'd42];

assign tmp_651_fu_17431_p3 = r_V_79_fu_484_p2[32'd23];

assign tmp_654_fu_19244_p3 = r_V_79_reg_9079[32'd43];

assign tmp_657_fu_17495_p3 = r_V_80_fu_509_p2[32'd23];

assign tmp_660_fu_19369_p3 = r_V_80_reg_9083[32'd41];

assign tmp_663_fu_17559_p3 = r_V_81_fu_489_p2[32'd23];

assign tmp_666_fu_19494_p3 = r_V_81_reg_9087[32'd41];

assign tmp_669_fu_17623_p3 = r_V_82_fu_497_p2[32'd23];

assign tmp_672_fu_19619_p3 = r_V_82_reg_9091[32'd43];

assign tmp_675_fu_17687_p3 = r_V_83_fu_507_p2[32'd23];

assign tmp_678_fu_19744_p3 = r_V_83_reg_9095[32'd44];

assign tmp_681_fu_17751_p3 = r_V_84_fu_494_p2[32'd23];

assign tmp_684_fu_19869_p3 = r_V_84_reg_9099[32'd39];

assign tmp_687_fu_17815_p3 = r_V_85_fu_495_p2[32'd23];

assign tmp_690_fu_19994_p3 = r_V_85_reg_9103[32'd42];

assign tmp_696_fu_20142_p3 = r_V_86_reg_9107[32'd44];

assign tmp_702_fu_20291_p3 = r_V_87_reg_9111[32'd41];

assign tmp_708_fu_20440_p3 = r_V_88_reg_9115[32'd39];

assign tmp_714_fu_20589_p3 = r_V_89_reg_9119[32'd43];

assign tmp_720_fu_20738_p3 = r_V_90_reg_9123[32'd41];

assign tmp_723_fu_18157_p3 = r_V_91_fu_18121_p2[32'd23];

assign tmp_726_fu_18221_p3 = r_V_91_fu_18121_p2[32'd39];

assign tmp_732_fu_20904_p3 = r_V_92_reg_9127[32'd41];

assign tmp_738_fu_21053_p3 = r_V_93_reg_9131[32'd42];

assign tmp_744_fu_21202_p3 = r_V_94_reg_9135[32'd38];

assign tmp_750_fu_21347_p3 = r_V_95_reg_9139[32'd54];

assign tmp_756_fu_21492_p3 = r_V_96_reg_9143[32'd43];

assign tmp_762_fu_21621_p3 = r_V_97_reg_9147[32'd40];

assign tmp_768_fu_21746_p3 = r_V_98_reg_9151[32'd55];

assign tmp_774_fu_21891_p3 = r_V_99_reg_9155[32'd51];

assign tmp_780_fu_22020_p3 = r_V_100_reg_9159[32'd44];

assign tmp_786_fu_22149_p3 = r_V_101_reg_9163[32'd42];

assign tmp_792_fu_22278_p3 = r_V_102_reg_9167[32'd40];

assign tmp_798_fu_22407_p3 = r_V_103_reg_9171[32'd46];

assign tmp_801_fu_22536_p3 = r_V_104_fu_466_p2[32'd23];

assign tmp_804_fu_25569_p3 = r_V_104_reg_12983[32'd41];

assign tmp_807_fu_22600_p3 = r_V_105_fu_539_p2[32'd23];

assign tmp_810_fu_25694_p3 = r_V_105_reg_12987[32'd42];

assign tmp_813_fu_22664_p3 = r_V_106_fu_512_p2[32'd23];

assign tmp_816_fu_25819_p3 = r_V_106_reg_12991[32'd41];

assign tmp_819_fu_22728_p3 = r_V_107_fu_463_p2[32'd23];

assign tmp_822_fu_25944_p3 = r_V_107_reg_12995[32'd42];

assign tmp_825_fu_22792_p3 = r_V_108_fu_529_p2[32'd23];

assign tmp_828_fu_26069_p3 = r_V_108_reg_12999[32'd43];

assign tmp_831_fu_22856_p3 = r_V_109_fu_485_p2[32'd23];

assign tmp_834_fu_26194_p3 = r_V_109_reg_13003[32'd41];

assign tmp_840_fu_23003_p3 = r_V_110_fu_22912_p2[32'd38];

assign tmp_843_fu_23119_p3 = r_V_111_fu_526_p2[32'd23];

assign tmp_846_fu_26336_p3 = r_V_111_reg_13007[32'd43];

assign tmp_849_fu_23183_p3 = r_V_112_fu_471_p2[32'd23];

assign tmp_852_fu_26461_p3 = r_V_112_reg_13011[32'd42];

assign tmp_858_fu_26605_p3 = r_V_113_reg_13015[32'd54];

assign tmp_864_fu_26754_p3 = r_V_114_reg_13019[32'd41];

assign tmp_870_fu_26903_p3 = r_V_115_reg_13023[32'd44];

assign tmp_876_fu_27052_p3 = r_V_116_reg_13027[32'd44];

assign tmp_882_fu_27201_p3 = r_V_117_reg_13031[32'd46];

assign tmp_888_fu_27350_p3 = r_V_118_reg_13035[32'd42];

assign tmp_894_fu_27499_p3 = r_V_119_reg_13039[32'd44];

assign tmp_900_fu_27648_p3 = r_V_120_reg_13043[32'd43];

assign tmp_906_fu_27797_p3 = r_V_121_reg_13047[32'd43];

assign tmp_912_fu_28031_p3 = r_V_122_fu_27940_p2[32'd40];

assign tmp_915_fu_28147_p3 = r_V_123_fu_472_p2[32'd23];

assign tmp_918_fu_31367_p3 = r_V_123_reg_15547[32'd42];

assign tmp_921_fu_28211_p3 = r_V_124_fu_462_p2[32'd23];

assign tmp_924_fu_31492_p3 = r_V_124_reg_15551[32'd43];

assign tmp_927_fu_28275_p3 = r_V_125_fu_510_p2[32'd23];

assign tmp_930_fu_31617_p3 = r_V_125_reg_15555[32'd42];

assign tmp_933_fu_28339_p3 = r_V_126_fu_515_p2[32'd23];

assign tmp_936_fu_31742_p3 = r_V_126_reg_15559[32'd43];

assign tmp_939_fu_28403_p3 = r_V_127_fu_479_p2[32'd23];

assign tmp_942_fu_31867_p3 = r_V_127_reg_15563[32'd42];

assign tmp_945_fu_28467_p3 = r_V_128_fu_513_p2[32'd23];

assign tmp_948_fu_31992_p3 = r_V_128_reg_15567[32'd44];

assign tmp_951_fu_28531_p3 = r_V_129_fu_521_p2[32'd23];

assign tmp_954_fu_32117_p3 = r_V_129_reg_15571[32'd39];

assign tmp_957_fu_28595_p3 = r_V_130_fu_491_p2[32'd23];

assign tmp_960_fu_32242_p3 = r_V_130_reg_15575[32'd41];

assign tmp_966_fu_32390_p3 = r_V_131_reg_15579[32'd43];

assign tmp_972_fu_32539_p3 = r_V_132_reg_15583[32'd42];

assign tmp_978_fu_32688_p3 = r_V_133_reg_15587[32'd42];

assign tmp_984_fu_32837_p3 = r_V_134_reg_15591[32'd43];

assign tmp_990_fu_32986_p3 = r_V_135_reg_15595[32'd42];

assign tmp_996_fu_33135_p3 = r_V_136_reg_15599[32'd42];

assign tmp_fu_17303_p3 = r_V_fu_536_p2[32'd23];

assign trunc_ln1273_10_fu_18928_p0 = p_read6_int_reg;

assign trunc_ln1273_10_fu_18928_p1 = trunc_ln1273_10_fu_18928_p0[15:0];

assign trunc_ln1273_11_fu_18940_p0 = p_read6_int_reg;

assign trunc_ln1273_11_fu_18940_p1 = trunc_ln1273_11_fu_18940_p0[18:0];

assign trunc_ln1273_2_fu_18868_p3 = {{trunc_ln1273_7_fu_18864_p1}, {1'd0}};

assign trunc_ln1273_3_fu_18894_p3 = {{trunc_ln1273_8_fu_18890_p1}, {8'd0}};

assign trunc_ln1273_4_fu_18906_p3 = {{trunc_ln1273_9_fu_18902_p1}, {1'd0}};

assign trunc_ln1273_5_fu_18932_p3 = {{trunc_ln1273_10_fu_18928_p1}, {8'd0}};

assign trunc_ln1273_6_fu_18944_p3 = {{trunc_ln1273_11_fu_18940_p1}, {5'd0}};

assign trunc_ln1273_7_fu_18864_p0 = p_read3_int_reg;

assign trunc_ln1273_7_fu_18864_p1 = trunc_ln1273_7_fu_18864_p0[22:0];

assign trunc_ln1273_8_fu_18890_p0 = p_read5_int_reg;

assign trunc_ln1273_8_fu_18890_p1 = trunc_ln1273_8_fu_18890_p0[15:0];

assign trunc_ln1273_9_fu_18902_p0 = p_read5_int_reg;

assign trunc_ln1273_9_fu_18902_p1 = trunc_ln1273_9_fu_18902_p0[22:0];

assign trunc_ln1273_fu_18852_p0 = p_read3_int_reg;

assign trunc_ln1273_fu_18852_p1 = trunc_ln1273_fu_18852_p0[17:0];

assign trunc_ln5_fu_18856_p3 = {{trunc_ln1273_fu_18852_p1}, {6'd0}};

assign underflow_162_fu_19189_p2 = (xor_ln896_486_fu_19183_p2 & p_Result_405_reg_41364);

assign underflow_163_fu_19314_p2 = (xor_ln896_487_fu_19308_p2 & p_Result_408_reg_41395);

assign underflow_164_fu_19439_p2 = (xor_ln896_488_fu_19433_p2 & p_Result_411_reg_41426);

assign underflow_165_fu_19564_p2 = (xor_ln896_489_fu_19558_p2 & p_Result_414_reg_41457);

assign underflow_166_fu_19689_p2 = (xor_ln896_490_fu_19683_p2 & p_Result_417_reg_41488);

assign underflow_167_fu_19814_p2 = (xor_ln896_491_fu_19808_p2 & p_Result_420_reg_41519);

assign underflow_168_fu_19939_p2 = (xor_ln896_492_fu_19933_p2 & p_Result_423_reg_41550);

assign underflow_169_fu_20064_p2 = (xor_ln896_493_fu_20058_p2 & p_Result_426_reg_41581);

assign underflow_170_fu_20213_p2 = (xor_ln896_494_fu_20207_p2 & p_Result_429_reg_41612);

assign underflow_171_fu_20362_p2 = (xor_ln896_495_fu_20356_p2 & p_Result_432_reg_41641);

assign underflow_172_fu_20511_p2 = (xor_ln896_496_fu_20505_p2 & p_Result_435_reg_41670);

assign underflow_173_fu_20660_p2 = (xor_ln896_497_fu_20654_p2 & p_Result_438_reg_41699);

assign underflow_174_fu_20809_p2 = (xor_ln896_498_fu_20803_p2 & p_Result_441_reg_41728);

assign underflow_175_fu_18295_p2 = (xor_ln896_499_fu_18289_p2 & p_Result_444_fu_18127_p3);

assign underflow_176_fu_20975_p2 = (xor_ln896_500_fu_20969_p2 & p_Result_447_reg_41772);

assign underflow_177_fu_21124_p2 = (xor_ln896_501_fu_21118_p2 & p_Result_450_reg_41801);

assign underflow_178_fu_21273_p2 = (xor_ln896_502_fu_21267_p2 & p_Result_453_reg_41830);

assign underflow_179_fu_21418_p2 = (xor_ln896_503_fu_21412_p2 & p_Result_456_reg_41859);

assign underflow_180_fu_21563_p2 = (xor_ln896_504_fu_21557_p2 & p_Result_459_reg_41888);

assign underflow_181_fu_21692_p2 = (xor_ln896_505_fu_21686_p2 & p_Result_462_reg_41917);

assign underflow_182_fu_21817_p2 = (xor_ln896_506_fu_21811_p2 & p_Result_465_reg_41946);

assign underflow_183_fu_21962_p2 = (xor_ln896_507_fu_21956_p2 & p_Result_468_reg_41975);

assign underflow_184_fu_22091_p2 = (xor_ln896_508_fu_22085_p2 & p_Result_471_reg_42004);

assign underflow_185_fu_22220_p2 = (xor_ln896_509_fu_22214_p2 & p_Result_474_reg_42033);

assign underflow_186_fu_22349_p2 = (xor_ln896_510_fu_22343_p2 & p_Result_477_reg_42062);

assign underflow_187_fu_22478_p2 = (xor_ln896_511_fu_22472_p2 & p_Result_480_reg_42091);

assign underflow_188_fu_25639_p2 = (xor_ln896_512_fu_25633_p2 & p_Result_483_reg_42252);

assign underflow_189_fu_25764_p2 = (xor_ln896_513_fu_25758_p2 & p_Result_486_reg_42283);

assign underflow_190_fu_25889_p2 = (xor_ln896_514_fu_25883_p2 & p_Result_489_reg_42314);

assign underflow_191_fu_26014_p2 = (xor_ln896_515_fu_26008_p2 & p_Result_492_reg_42345);

assign underflow_192_fu_26139_p2 = (xor_ln896_516_fu_26133_p2 & p_Result_495_reg_42376);

assign underflow_193_fu_26264_p2 = (xor_ln896_517_fu_26258_p2 & p_Result_498_reg_42407);

assign underflow_194_fu_23077_p2 = (xor_ln896_518_fu_23071_p2 & p_Result_501_fu_22918_p3);

assign underflow_195_fu_26406_p2 = (xor_ln896_519_fu_26400_p2 & p_Result_504_reg_42453);

assign underflow_196_fu_26531_p2 = (xor_ln896_520_fu_26525_p2 & p_Result_507_reg_42484);

assign underflow_197_fu_26676_p2 = (xor_ln896_521_fu_26670_p2 & p_Result_510_reg_42515);

assign underflow_198_fu_26825_p2 = (xor_ln896_522_fu_26819_p2 & p_Result_513_reg_42544);

assign underflow_199_fu_26974_p2 = (xor_ln896_523_fu_26968_p2 & p_Result_516_reg_42573);

assign underflow_200_fu_27123_p2 = (xor_ln896_524_fu_27117_p2 & p_Result_519_reg_42602);

assign underflow_201_fu_27272_p2 = (xor_ln896_525_fu_27266_p2 & p_Result_522_reg_42631);

assign underflow_202_fu_27421_p2 = (xor_ln896_526_fu_27415_p2 & p_Result_525_reg_42660);

assign underflow_203_fu_27570_p2 = (xor_ln896_527_fu_27564_p2 & p_Result_528_reg_42689);

assign underflow_204_fu_27719_p2 = (xor_ln896_528_fu_27713_p2 & p_Result_531_reg_42718);

assign underflow_205_fu_27868_p2 = (xor_ln896_529_fu_27862_p2 & p_Result_534_reg_42747);

assign underflow_206_fu_28105_p2 = (xor_ln896_530_fu_28099_p2 & p_Result_537_fu_27946_p3);

assign underflow_207_fu_31437_p2 = (xor_ln896_531_fu_31431_p2 & p_Result_540_reg_42845);

assign underflow_208_fu_31562_p2 = (xor_ln896_532_fu_31556_p2 & p_Result_543_reg_42876);

assign underflow_209_fu_31687_p2 = (xor_ln896_533_fu_31681_p2 & p_Result_546_reg_42907);

assign underflow_210_fu_31812_p2 = (xor_ln896_534_fu_31806_p2 & p_Result_549_reg_42938);

assign underflow_211_fu_31937_p2 = (xor_ln896_535_fu_31931_p2 & p_Result_552_reg_42969);

assign underflow_212_fu_32062_p2 = (xor_ln896_536_fu_32056_p2 & p_Result_555_reg_43000);

assign underflow_213_fu_32187_p2 = (xor_ln896_537_fu_32181_p2 & p_Result_558_reg_43031);

assign underflow_214_fu_32312_p2 = (xor_ln896_538_fu_32306_p2 & p_Result_561_reg_43062);

assign underflow_215_fu_32461_p2 = (xor_ln896_539_fu_32455_p2 & p_Result_564_reg_43093);

assign underflow_216_fu_32610_p2 = (xor_ln896_540_fu_32604_p2 & p_Result_567_reg_43122);

assign underflow_217_fu_32759_p2 = (xor_ln896_541_fu_32753_p2 & p_Result_570_reg_43151);

assign underflow_218_fu_32908_p2 = (xor_ln896_542_fu_32902_p2 & p_Result_573_reg_43180);

assign underflow_219_fu_33057_p2 = (xor_ln896_543_fu_33051_p2 & p_Result_576_reg_43209);

assign underflow_220_fu_33206_p2 = (xor_ln896_544_fu_33200_p2 & p_Result_579_reg_43238);

assign underflow_221_fu_33355_p2 = (xor_ln896_545_fu_33349_p2 & p_Result_582_reg_43267);

assign underflow_222_fu_33504_p2 = (xor_ln896_546_fu_33498_p2 & p_Result_585_reg_43296);

assign underflow_223_fu_29172_p2 = (xor_ln896_547_fu_29166_p2 & p_Result_588_fu_29013_p3);

assign underflow_224_fu_37171_p2 = (xor_ln896_548_fu_37165_p2 & p_Result_591_reg_43520);

assign underflow_225_fu_37295_p2 = (xor_ln896_549_fu_37289_p2 & p_Result_594_reg_43551);

assign underflow_226_fu_37420_p2 = (xor_ln896_550_fu_37414_p2 & p_Result_597_reg_43582);

assign underflow_227_fu_37545_p2 = (xor_ln896_551_fu_37539_p2 & p_Result_600_reg_43613);

assign underflow_228_fu_37670_p2 = (xor_ln896_552_fu_37664_p2 & p_Result_603_reg_43644);

assign underflow_229_fu_37795_p2 = (xor_ln896_553_fu_37789_p2 & p_Result_606_reg_43675);

assign underflow_230_fu_37920_p2 = (xor_ln896_554_fu_37914_p2 & p_Result_609_reg_43706);

assign underflow_231_fu_38045_p2 = (xor_ln896_555_fu_38039_p2 & p_Result_612_reg_43737);

assign underflow_232_fu_38170_p2 = (xor_ln896_556_fu_38164_p2 & p_Result_615_reg_43768);

assign underflow_233_fu_38315_p2 = (xor_ln896_557_fu_38309_p2 & p_Result_618_reg_43799);

assign underflow_234_fu_38464_p2 = (xor_ln896_558_fu_38458_p2 & p_Result_621_reg_43828);

assign underflow_235_fu_38613_p2 = (xor_ln896_559_fu_38607_p2 & p_Result_624_reg_43857);

assign underflow_236_fu_38762_p2 = (xor_ln896_560_fu_38756_p2 & p_Result_627_reg_43886);

assign underflow_237_fu_38911_p2 = (xor_ln896_561_fu_38905_p2 & p_Result_630_reg_43915);

assign underflow_238_fu_39060_p2 = (xor_ln896_562_fu_39054_p2 & p_Result_633_reg_43944);

assign underflow_239_fu_39209_p2 = (xor_ln896_563_fu_39203_p2 & p_Result_636_reg_43973);

assign underflow_240_fu_34664_p2 = (xor_ln896_564_fu_34658_p2 & p_Result_639_fu_34496_p3);

assign underflow_241_fu_39375_p2 = (xor_ln896_565_fu_39369_p2 & p_Result_642_reg_44017);

assign underflow_242_fu_23672_p2 = (xor_ln896_404_fu_23666_p2 & p_Result_645_fu_23632_p3);

assign underflow_243_fu_23770_p2 = (xor_ln896_405_fu_23764_p2 & p_Result_647_fu_23730_p3);

assign underflow_244_fu_23868_p2 = (xor_ln896_406_fu_23862_p2 & p_Result_649_fu_23828_p3);

assign underflow_245_fu_23966_p2 = (xor_ln896_407_fu_23960_p2 & p_Result_651_fu_23926_p3);

assign underflow_246_fu_24064_p2 = (xor_ln896_408_fu_24058_p2 & p_Result_653_fu_24024_p3);

assign underflow_247_fu_24162_p2 = (xor_ln896_409_fu_24156_p2 & p_Result_655_fu_24122_p3);

assign underflow_248_fu_24260_p2 = (xor_ln896_410_fu_24254_p2 & p_Result_657_fu_24220_p3);

assign underflow_249_fu_24358_p2 = (xor_ln896_411_fu_24352_p2 & p_Result_659_fu_24318_p3);

assign underflow_250_fu_24456_p2 = (xor_ln896_412_fu_24450_p2 & p_Result_661_fu_24416_p3);

assign underflow_251_fu_24558_p2 = (xor_ln896_413_fu_24552_p2 & p_Result_663_fu_24518_p3);

assign underflow_252_fu_24660_p2 = (xor_ln896_414_fu_24654_p2 & p_Result_665_fu_24620_p3);

assign underflow_253_fu_24762_p2 = (xor_ln896_415_fu_24756_p2 & p_Result_667_fu_24722_p3);

assign underflow_254_fu_24864_p2 = (xor_ln896_416_fu_24858_p2 & p_Result_669_fu_24824_p3);

assign underflow_255_fu_24966_p2 = (xor_ln896_417_fu_24960_p2 & p_Result_671_fu_24926_p3);

assign underflow_256_fu_25068_p2 = (xor_ln896_418_fu_25062_p2 & p_Result_673_fu_25028_p3);

assign underflow_257_fu_25170_p2 = (xor_ln896_419_fu_25164_p2 & p_Result_675_fu_25130_p3);

assign underflow_258_fu_25272_p2 = (xor_ln896_420_fu_25266_p2 & p_Result_677_fu_25232_p3);

assign underflow_259_fu_25374_p2 = (xor_ln896_421_fu_25368_p2 & p_Result_679_fu_25334_p3);

assign underflow_260_fu_29234_p2 = (xor_ln896_422_fu_29228_p2 & p_Result_681_fu_29196_p3);

assign underflow_261_fu_29334_p2 = (xor_ln896_423_fu_29328_p2 & p_Result_683_fu_29295_p3);

assign underflow_262_fu_29434_p2 = (xor_ln896_424_fu_29428_p2 & p_Result_685_fu_29395_p3);

assign underflow_263_fu_29532_p2 = (xor_ln896_425_fu_29526_p2 & p_Result_687_fu_29494_p3);

assign underflow_264_fu_29632_p2 = (xor_ln896_426_fu_29626_p2 & p_Result_689_fu_29593_p3);

assign underflow_265_fu_29732_p2 = (xor_ln896_427_fu_29726_p2 & p_Result_691_fu_29693_p3);

assign underflow_266_fu_29832_p2 = (xor_ln896_428_fu_29826_p2 & p_Result_693_fu_29793_p3);

assign underflow_267_fu_29932_p2 = (xor_ln896_429_fu_29926_p2 & p_Result_695_fu_29893_p3);

assign underflow_268_fu_30032_p2 = (xor_ln896_430_fu_30026_p2 & p_Result_697_fu_29993_p3);

assign underflow_269_fu_30134_p2 = (xor_ln896_431_fu_30128_p2 & p_Result_699_fu_30094_p3);

assign underflow_270_fu_30236_p2 = (xor_ln896_432_fu_30230_p2 & p_Result_701_fu_30196_p3);

assign underflow_271_fu_30338_p2 = (xor_ln896_433_fu_30332_p2 & p_Result_703_fu_30298_p3);

assign underflow_272_fu_30440_p2 = (xor_ln896_434_fu_30434_p2 & p_Result_705_fu_30400_p3);

assign underflow_273_fu_30542_p2 = (xor_ln896_435_fu_30536_p2 & p_Result_707_fu_30502_p3);

assign underflow_274_fu_30644_p2 = (xor_ln896_436_fu_30638_p2 & p_Result_709_fu_30604_p3);

assign underflow_275_fu_30746_p2 = (xor_ln896_437_fu_30740_p2 & p_Result_711_fu_30706_p3);

assign underflow_276_fu_30848_p2 = (xor_ln896_438_fu_30842_p2 & p_Result_713_fu_30808_p3);

assign underflow_277_fu_30950_p2 = (xor_ln896_439_fu_30944_p2 & p_Result_715_fu_30910_p3);

assign underflow_278_fu_34733_p2 = (xor_ln896_440_fu_34728_p2 & p_Result_717_reg_43340);

assign underflow_279_fu_34791_p2 = (xor_ln896_441_fu_34786_p2 & p_Result_719_reg_43360);

assign underflow_280_fu_34849_p2 = (xor_ln896_442_fu_34844_p2 & p_Result_721_reg_43380);

assign underflow_281_fu_34907_p2 = (xor_ln896_443_fu_34902_p2 & p_Result_723_reg_43400);

assign underflow_282_fu_34965_p2 = (xor_ln896_444_fu_34960_p2 & p_Result_725_reg_43420);

assign underflow_283_fu_35023_p2 = (xor_ln896_445_fu_35018_p2 & p_Result_727_reg_43440);

assign underflow_284_fu_35081_p2 = (xor_ln896_446_fu_35076_p2 & p_Result_729_reg_43460);

assign underflow_285_fu_35139_p2 = (xor_ln896_447_fu_35134_p2 & p_Result_731_reg_43480);

assign underflow_286_fu_35197_p2 = (xor_ln896_448_fu_35192_p2 & p_Result_733_reg_43500);

assign underflow_287_fu_35294_p2 = (xor_ln896_449_fu_35288_p2 & p_Result_735_fu_35254_p3);

assign underflow_288_fu_35396_p2 = (xor_ln896_450_fu_35390_p2 & p_Result_737_fu_35356_p3);

assign underflow_289_fu_35498_p2 = (xor_ln896_451_fu_35492_p2 & p_Result_739_fu_35458_p3);

assign underflow_290_fu_35600_p2 = (xor_ln896_452_fu_35594_p2 & p_Result_741_fu_35560_p3);

assign underflow_291_fu_35702_p2 = (xor_ln896_453_fu_35696_p2 & p_Result_743_fu_35662_p3);

assign underflow_292_fu_35804_p2 = (xor_ln896_454_fu_35798_p2 & p_Result_745_fu_35764_p3);

assign underflow_293_fu_35906_p2 = (xor_ln896_455_fu_35900_p2 & p_Result_747_fu_35866_p3);

assign underflow_294_fu_36008_p2 = (xor_ln896_456_fu_36002_p2 & p_Result_749_fu_35968_p3);

assign underflow_295_fu_36110_p2 = (xor_ln896_457_fu_36104_p2 & p_Result_751_fu_36070_p3);

assign underflow_296_fu_36212_p2 = (xor_ln896_458_fu_36206_p2 & p_Result_753_fu_36172_p3);

assign underflow_297_fu_36314_p2 = (xor_ln896_459_fu_36308_p2 & p_Result_755_fu_36274_p3);

assign underflow_298_fu_36416_p2 = (xor_ln896_460_fu_36410_p2 & p_Result_757_fu_36376_p3);

assign underflow_299_fu_36518_p2 = (xor_ln896_461_fu_36512_p2 & p_Result_759_fu_36478_p3);

assign underflow_300_fu_36620_p2 = (xor_ln896_462_fu_36614_p2 & p_Result_761_fu_36580_p3);

assign underflow_301_fu_36722_p2 = (xor_ln896_463_fu_36716_p2 & p_Result_763_fu_36682_p3);

assign underflow_302_fu_36824_p2 = (xor_ln896_464_fu_36818_p2 & p_Result_765_fu_36784_p3);

assign underflow_303_fu_36926_p2 = (xor_ln896_465_fu_36920_p2 & p_Result_767_fu_36886_p3);

assign underflow_304_fu_37028_p2 = (xor_ln896_466_fu_37022_p2 & p_Result_769_fu_36988_p3);

assign underflow_305_fu_39454_p2 = (xor_ln896_467_fu_39448_p2 & p_Result_771_fu_39415_p3);

assign underflow_306_fu_39554_p2 = (xor_ln896_468_fu_39548_p2 & p_Result_773_fu_39515_p3);

assign underflow_307_fu_39654_p2 = (xor_ln896_469_fu_39648_p2 & p_Result_775_fu_39615_p3);

assign underflow_308_fu_39754_p2 = (xor_ln896_470_fu_39748_p2 & p_Result_777_fu_39715_p3);

assign underflow_309_fu_39854_p2 = (xor_ln896_471_fu_39848_p2 & p_Result_779_fu_39815_p3);

assign underflow_310_fu_39954_p2 = (xor_ln896_472_fu_39948_p2 & p_Result_781_fu_39915_p3);

assign underflow_311_fu_40054_p2 = (xor_ln896_473_fu_40048_p2 & p_Result_783_fu_40015_p3);

assign underflow_312_fu_40154_p2 = (xor_ln896_474_fu_40148_p2 & p_Result_785_fu_40115_p3);

assign underflow_313_fu_40254_p2 = (xor_ln896_475_fu_40248_p2 & p_Result_787_fu_40215_p3);

assign underflow_314_fu_40356_p2 = (xor_ln896_476_fu_40350_p2 & p_Result_789_fu_40316_p3);

assign underflow_315_fu_40458_p2 = (xor_ln896_477_fu_40452_p2 & p_Result_791_fu_40418_p3);

assign underflow_316_fu_40560_p2 = (xor_ln896_478_fu_40554_p2 & p_Result_793_fu_40520_p3);

assign underflow_317_fu_40662_p2 = (xor_ln896_479_fu_40656_p2 & p_Result_795_fu_40622_p3);

assign underflow_318_fu_40764_p2 = (xor_ln896_480_fu_40758_p2 & p_Result_797_fu_40724_p3);

assign underflow_319_fu_40866_p2 = (xor_ln896_481_fu_40860_p2 & p_Result_799_fu_40826_p3);

assign underflow_320_fu_40968_p2 = (xor_ln896_482_fu_40962_p2 & p_Result_801_fu_40928_p3);

assign underflow_321_fu_41070_p2 = (xor_ln896_483_fu_41064_p2 & p_Result_803_fu_41030_p3);

assign underflow_322_fu_41172_p2 = (xor_ln896_484_fu_41166_p2 & p_Result_805_fu_41132_p3);

assign underflow_fu_19064_p2 = (xor_ln896_485_fu_19058_p2 & p_Result_s_reg_41333);

assign xor_ln302_162_fu_23684_p2 = (xor_ln302_fu_23678_p2 ^ 1'd1);

assign xor_ln302_163_fu_23776_p2 = (p_Result_648_fu_23744_p3 ^ p_Result_647_fu_23730_p3);

assign xor_ln302_164_fu_23782_p2 = (xor_ln302_163_fu_23776_p2 ^ 1'd1);

assign xor_ln302_165_fu_23874_p2 = (p_Result_650_fu_23842_p3 ^ p_Result_649_fu_23828_p3);

assign xor_ln302_166_fu_23880_p2 = (xor_ln302_165_fu_23874_p2 ^ 1'd1);

assign xor_ln302_167_fu_23972_p2 = (p_Result_652_fu_23940_p3 ^ p_Result_651_fu_23926_p3);

assign xor_ln302_168_fu_23978_p2 = (xor_ln302_167_fu_23972_p2 ^ 1'd1);

assign xor_ln302_169_fu_24070_p2 = (p_Result_654_fu_24038_p3 ^ p_Result_653_fu_24024_p3);

assign xor_ln302_170_fu_24076_p2 = (xor_ln302_169_fu_24070_p2 ^ 1'd1);

assign xor_ln302_171_fu_24168_p2 = (p_Result_656_fu_24136_p3 ^ p_Result_655_fu_24122_p3);

assign xor_ln302_172_fu_24174_p2 = (xor_ln302_171_fu_24168_p2 ^ 1'd1);

assign xor_ln302_173_fu_24266_p2 = (p_Result_658_fu_24234_p3 ^ p_Result_657_fu_24220_p3);

assign xor_ln302_174_fu_24272_p2 = (xor_ln302_173_fu_24266_p2 ^ 1'd1);

assign xor_ln302_175_fu_24364_p2 = (p_Result_660_fu_24332_p3 ^ p_Result_659_fu_24318_p3);

assign xor_ln302_176_fu_24370_p2 = (xor_ln302_175_fu_24364_p2 ^ 1'd1);

assign xor_ln302_177_fu_24462_p2 = (p_Result_662_fu_24430_p3 ^ p_Result_661_fu_24416_p3);

assign xor_ln302_178_fu_24468_p2 = (xor_ln302_177_fu_24462_p2 ^ 1'd1);

assign xor_ln302_179_fu_24564_p2 = (p_Result_664_fu_24532_p3 ^ p_Result_663_fu_24518_p3);

assign xor_ln302_180_fu_24570_p2 = (xor_ln302_179_fu_24564_p2 ^ 1'd1);

assign xor_ln302_181_fu_24666_p2 = (p_Result_666_fu_24634_p3 ^ p_Result_665_fu_24620_p3);

assign xor_ln302_182_fu_24672_p2 = (xor_ln302_181_fu_24666_p2 ^ 1'd1);

assign xor_ln302_183_fu_24768_p2 = (p_Result_668_fu_24736_p3 ^ p_Result_667_fu_24722_p3);

assign xor_ln302_184_fu_24774_p2 = (xor_ln302_183_fu_24768_p2 ^ 1'd1);

assign xor_ln302_185_fu_24870_p2 = (p_Result_670_fu_24838_p3 ^ p_Result_669_fu_24824_p3);

assign xor_ln302_186_fu_24876_p2 = (xor_ln302_185_fu_24870_p2 ^ 1'd1);

assign xor_ln302_187_fu_24972_p2 = (p_Result_672_fu_24940_p3 ^ p_Result_671_fu_24926_p3);

assign xor_ln302_188_fu_24978_p2 = (xor_ln302_187_fu_24972_p2 ^ 1'd1);

assign xor_ln302_189_fu_25074_p2 = (p_Result_674_fu_25042_p3 ^ p_Result_673_fu_25028_p3);

assign xor_ln302_190_fu_25080_p2 = (xor_ln302_189_fu_25074_p2 ^ 1'd1);

assign xor_ln302_191_fu_25176_p2 = (p_Result_676_fu_25144_p3 ^ p_Result_675_fu_25130_p3);

assign xor_ln302_192_fu_25182_p2 = (xor_ln302_191_fu_25176_p2 ^ 1'd1);

assign xor_ln302_193_fu_25278_p2 = (p_Result_678_fu_25246_p3 ^ p_Result_677_fu_25232_p3);

assign xor_ln302_194_fu_25284_p2 = (xor_ln302_193_fu_25278_p2 ^ 1'd1);

assign xor_ln302_195_fu_25380_p2 = (p_Result_680_fu_25348_p3 ^ p_Result_679_fu_25334_p3);

assign xor_ln302_196_fu_25386_p2 = (xor_ln302_195_fu_25380_p2 ^ 1'd1);

assign xor_ln302_197_fu_29240_p2 = (p_Result_682_fu_29208_p3 ^ p_Result_681_fu_29196_p3);

assign xor_ln302_198_fu_29246_p2 = (xor_ln302_197_fu_29240_p2 ^ 1'd1);

assign xor_ln302_199_fu_29340_p2 = (p_Result_684_fu_29308_p3 ^ p_Result_683_fu_29295_p3);

assign xor_ln302_200_fu_29346_p2 = (xor_ln302_199_fu_29340_p2 ^ 1'd1);

assign xor_ln302_201_fu_29440_p2 = (p_Result_686_fu_29408_p3 ^ p_Result_685_fu_29395_p3);

assign xor_ln302_202_fu_29446_p2 = (xor_ln302_201_fu_29440_p2 ^ 1'd1);

assign xor_ln302_203_fu_29538_p2 = (p_Result_688_fu_29506_p3 ^ p_Result_687_fu_29494_p3);

assign xor_ln302_204_fu_29544_p2 = (xor_ln302_203_fu_29538_p2 ^ 1'd1);

assign xor_ln302_205_fu_29638_p2 = (p_Result_690_fu_29606_p3 ^ p_Result_689_fu_29593_p3);

assign xor_ln302_206_fu_29644_p2 = (xor_ln302_205_fu_29638_p2 ^ 1'd1);

assign xor_ln302_207_fu_29738_p2 = (p_Result_692_fu_29706_p3 ^ p_Result_691_fu_29693_p3);

assign xor_ln302_208_fu_29744_p2 = (xor_ln302_207_fu_29738_p2 ^ 1'd1);

assign xor_ln302_209_fu_29838_p2 = (p_Result_694_fu_29806_p3 ^ p_Result_693_fu_29793_p3);

assign xor_ln302_210_fu_29844_p2 = (xor_ln302_209_fu_29838_p2 ^ 1'd1);

assign xor_ln302_211_fu_29938_p2 = (p_Result_696_fu_29906_p3 ^ p_Result_695_fu_29893_p3);

assign xor_ln302_212_fu_29944_p2 = (xor_ln302_211_fu_29938_p2 ^ 1'd1);

assign xor_ln302_213_fu_30038_p2 = (p_Result_698_fu_30006_p3 ^ p_Result_697_fu_29993_p3);

assign xor_ln302_214_fu_30044_p2 = (xor_ln302_213_fu_30038_p2 ^ 1'd1);

assign xor_ln302_215_fu_30140_p2 = (p_Result_700_fu_30108_p3 ^ p_Result_699_fu_30094_p3);

assign xor_ln302_216_fu_30146_p2 = (xor_ln302_215_fu_30140_p2 ^ 1'd1);

assign xor_ln302_217_fu_30242_p2 = (p_Result_702_fu_30210_p3 ^ p_Result_701_fu_30196_p3);

assign xor_ln302_218_fu_30248_p2 = (xor_ln302_217_fu_30242_p2 ^ 1'd1);

assign xor_ln302_219_fu_30344_p2 = (p_Result_704_fu_30312_p3 ^ p_Result_703_fu_30298_p3);

assign xor_ln302_220_fu_30350_p2 = (xor_ln302_219_fu_30344_p2 ^ 1'd1);

assign xor_ln302_221_fu_30446_p2 = (p_Result_706_fu_30414_p3 ^ p_Result_705_fu_30400_p3);

assign xor_ln302_222_fu_30452_p2 = (xor_ln302_221_fu_30446_p2 ^ 1'd1);

assign xor_ln302_223_fu_30548_p2 = (p_Result_708_fu_30516_p3 ^ p_Result_707_fu_30502_p3);

assign xor_ln302_224_fu_30554_p2 = (xor_ln302_223_fu_30548_p2 ^ 1'd1);

assign xor_ln302_225_fu_30650_p2 = (p_Result_710_fu_30618_p3 ^ p_Result_709_fu_30604_p3);

assign xor_ln302_226_fu_30656_p2 = (xor_ln302_225_fu_30650_p2 ^ 1'd1);

assign xor_ln302_227_fu_30752_p2 = (p_Result_712_fu_30720_p3 ^ p_Result_711_fu_30706_p3);

assign xor_ln302_228_fu_30758_p2 = (xor_ln302_227_fu_30752_p2 ^ 1'd1);

assign xor_ln302_229_fu_30854_p2 = (p_Result_714_fu_30822_p3 ^ p_Result_713_fu_30808_p3);

assign xor_ln302_230_fu_30860_p2 = (xor_ln302_229_fu_30854_p2 ^ 1'd1);

assign xor_ln302_231_fu_30956_p2 = (p_Result_716_fu_30924_p3 ^ p_Result_715_fu_30910_p3);

assign xor_ln302_232_fu_30962_p2 = (xor_ln302_231_fu_30956_p2 ^ 1'd1);

assign xor_ln302_233_fu_34738_p2 = (p_Result_718_reg_43353 ^ p_Result_717_reg_43340);

assign xor_ln302_234_fu_34742_p2 = (xor_ln302_233_fu_34738_p2 ^ 1'd1);

assign xor_ln302_235_fu_34796_p2 = (p_Result_720_reg_43373 ^ p_Result_719_reg_43360);

assign xor_ln302_236_fu_34800_p2 = (xor_ln302_235_fu_34796_p2 ^ 1'd1);

assign xor_ln302_237_fu_34854_p2 = (p_Result_722_reg_43393 ^ p_Result_721_reg_43380);

assign xor_ln302_238_fu_34858_p2 = (xor_ln302_237_fu_34854_p2 ^ 1'd1);

assign xor_ln302_239_fu_34912_p2 = (p_Result_724_reg_43413 ^ p_Result_723_reg_43400);

assign xor_ln302_240_fu_34916_p2 = (xor_ln302_239_fu_34912_p2 ^ 1'd1);

assign xor_ln302_241_fu_34970_p2 = (p_Result_726_reg_43433 ^ p_Result_725_reg_43420);

assign xor_ln302_242_fu_34974_p2 = (xor_ln302_241_fu_34970_p2 ^ 1'd1);

assign xor_ln302_243_fu_35028_p2 = (p_Result_728_reg_43453 ^ p_Result_727_reg_43440);

assign xor_ln302_244_fu_35032_p2 = (xor_ln302_243_fu_35028_p2 ^ 1'd1);

assign xor_ln302_245_fu_35086_p2 = (p_Result_730_reg_43473 ^ p_Result_729_reg_43460);

assign xor_ln302_246_fu_35090_p2 = (xor_ln302_245_fu_35086_p2 ^ 1'd1);

assign xor_ln302_247_fu_35144_p2 = (p_Result_732_reg_43493 ^ p_Result_731_reg_43480);

assign xor_ln302_248_fu_35148_p2 = (xor_ln302_247_fu_35144_p2 ^ 1'd1);

assign xor_ln302_249_fu_35202_p2 = (p_Result_734_reg_43513 ^ p_Result_733_reg_43500);

assign xor_ln302_250_fu_35206_p2 = (xor_ln302_249_fu_35202_p2 ^ 1'd1);

assign xor_ln302_251_fu_35300_p2 = (p_Result_736_fu_35268_p3 ^ p_Result_735_fu_35254_p3);

assign xor_ln302_252_fu_35306_p2 = (xor_ln302_251_fu_35300_p2 ^ 1'd1);

assign xor_ln302_253_fu_35402_p2 = (p_Result_738_fu_35370_p3 ^ p_Result_737_fu_35356_p3);

assign xor_ln302_254_fu_35408_p2 = (xor_ln302_253_fu_35402_p2 ^ 1'd1);

assign xor_ln302_255_fu_35504_p2 = (p_Result_740_fu_35472_p3 ^ p_Result_739_fu_35458_p3);

assign xor_ln302_256_fu_35510_p2 = (xor_ln302_255_fu_35504_p2 ^ 1'd1);

assign xor_ln302_257_fu_35606_p2 = (p_Result_742_fu_35574_p3 ^ p_Result_741_fu_35560_p3);

assign xor_ln302_258_fu_35612_p2 = (xor_ln302_257_fu_35606_p2 ^ 1'd1);

assign xor_ln302_259_fu_35708_p2 = (p_Result_744_fu_35676_p3 ^ p_Result_743_fu_35662_p3);

assign xor_ln302_260_fu_35714_p2 = (xor_ln302_259_fu_35708_p2 ^ 1'd1);

assign xor_ln302_261_fu_35810_p2 = (p_Result_746_fu_35778_p3 ^ p_Result_745_fu_35764_p3);

assign xor_ln302_262_fu_35816_p2 = (xor_ln302_261_fu_35810_p2 ^ 1'd1);

assign xor_ln302_263_fu_35912_p2 = (p_Result_748_fu_35880_p3 ^ p_Result_747_fu_35866_p3);

assign xor_ln302_264_fu_35918_p2 = (xor_ln302_263_fu_35912_p2 ^ 1'd1);

assign xor_ln302_265_fu_36014_p2 = (p_Result_750_fu_35982_p3 ^ p_Result_749_fu_35968_p3);

assign xor_ln302_266_fu_36020_p2 = (xor_ln302_265_fu_36014_p2 ^ 1'd1);

assign xor_ln302_267_fu_36116_p2 = (p_Result_752_fu_36084_p3 ^ p_Result_751_fu_36070_p3);

assign xor_ln302_268_fu_36122_p2 = (xor_ln302_267_fu_36116_p2 ^ 1'd1);

assign xor_ln302_269_fu_36218_p2 = (p_Result_754_fu_36186_p3 ^ p_Result_753_fu_36172_p3);

assign xor_ln302_270_fu_36224_p2 = (xor_ln302_269_fu_36218_p2 ^ 1'd1);

assign xor_ln302_271_fu_36320_p2 = (p_Result_756_fu_36288_p3 ^ p_Result_755_fu_36274_p3);

assign xor_ln302_272_fu_36326_p2 = (xor_ln302_271_fu_36320_p2 ^ 1'd1);

assign xor_ln302_273_fu_36422_p2 = (p_Result_758_fu_36390_p3 ^ p_Result_757_fu_36376_p3);

assign xor_ln302_274_fu_36428_p2 = (xor_ln302_273_fu_36422_p2 ^ 1'd1);

assign xor_ln302_275_fu_36524_p2 = (p_Result_760_fu_36492_p3 ^ p_Result_759_fu_36478_p3);

assign xor_ln302_276_fu_36530_p2 = (xor_ln302_275_fu_36524_p2 ^ 1'd1);

assign xor_ln302_277_fu_36626_p2 = (p_Result_762_fu_36594_p3 ^ p_Result_761_fu_36580_p3);

assign xor_ln302_278_fu_36632_p2 = (xor_ln302_277_fu_36626_p2 ^ 1'd1);

assign xor_ln302_279_fu_36728_p2 = (p_Result_764_fu_36696_p3 ^ p_Result_763_fu_36682_p3);

assign xor_ln302_280_fu_36734_p2 = (xor_ln302_279_fu_36728_p2 ^ 1'd1);

assign xor_ln302_281_fu_36830_p2 = (p_Result_766_fu_36798_p3 ^ p_Result_765_fu_36784_p3);

assign xor_ln302_282_fu_36836_p2 = (xor_ln302_281_fu_36830_p2 ^ 1'd1);

assign xor_ln302_283_fu_36932_p2 = (p_Result_768_fu_36900_p3 ^ p_Result_767_fu_36886_p3);

assign xor_ln302_284_fu_36938_p2 = (xor_ln302_283_fu_36932_p2 ^ 1'd1);

assign xor_ln302_285_fu_37034_p2 = (p_Result_770_fu_37002_p3 ^ p_Result_769_fu_36988_p3);

assign xor_ln302_286_fu_37040_p2 = (xor_ln302_285_fu_37034_p2 ^ 1'd1);

assign xor_ln302_287_fu_39460_p2 = (p_Result_772_fu_39428_p3 ^ p_Result_771_fu_39415_p3);

assign xor_ln302_288_fu_39466_p2 = (xor_ln302_287_fu_39460_p2 ^ 1'd1);

assign xor_ln302_289_fu_39560_p2 = (p_Result_774_fu_39528_p3 ^ p_Result_773_fu_39515_p3);

assign xor_ln302_290_fu_39566_p2 = (xor_ln302_289_fu_39560_p2 ^ 1'd1);

assign xor_ln302_291_fu_39660_p2 = (p_Result_776_fu_39628_p3 ^ p_Result_775_fu_39615_p3);

assign xor_ln302_292_fu_39666_p2 = (xor_ln302_291_fu_39660_p2 ^ 1'd1);

assign xor_ln302_293_fu_39760_p2 = (p_Result_778_fu_39728_p3 ^ p_Result_777_fu_39715_p3);

assign xor_ln302_294_fu_39766_p2 = (xor_ln302_293_fu_39760_p2 ^ 1'd1);

assign xor_ln302_295_fu_39860_p2 = (p_Result_780_fu_39828_p3 ^ p_Result_779_fu_39815_p3);

assign xor_ln302_296_fu_39866_p2 = (xor_ln302_295_fu_39860_p2 ^ 1'd1);

assign xor_ln302_297_fu_39960_p2 = (p_Result_782_fu_39928_p3 ^ p_Result_781_fu_39915_p3);

assign xor_ln302_298_fu_39966_p2 = (xor_ln302_297_fu_39960_p2 ^ 1'd1);

assign xor_ln302_299_fu_40060_p2 = (p_Result_784_fu_40028_p3 ^ p_Result_783_fu_40015_p3);

assign xor_ln302_300_fu_40066_p2 = (xor_ln302_299_fu_40060_p2 ^ 1'd1);

assign xor_ln302_301_fu_40160_p2 = (p_Result_786_fu_40128_p3 ^ p_Result_785_fu_40115_p3);

assign xor_ln302_302_fu_40166_p2 = (xor_ln302_301_fu_40160_p2 ^ 1'd1);

assign xor_ln302_303_fu_40260_p2 = (p_Result_788_fu_40228_p3 ^ p_Result_787_fu_40215_p3);

assign xor_ln302_304_fu_40266_p2 = (xor_ln302_303_fu_40260_p2 ^ 1'd1);

assign xor_ln302_305_fu_40362_p2 = (p_Result_790_fu_40330_p3 ^ p_Result_789_fu_40316_p3);

assign xor_ln302_306_fu_40368_p2 = (xor_ln302_305_fu_40362_p2 ^ 1'd1);

assign xor_ln302_307_fu_40464_p2 = (p_Result_792_fu_40432_p3 ^ p_Result_791_fu_40418_p3);

assign xor_ln302_308_fu_40470_p2 = (xor_ln302_307_fu_40464_p2 ^ 1'd1);

assign xor_ln302_309_fu_40566_p2 = (p_Result_794_fu_40534_p3 ^ p_Result_793_fu_40520_p3);

assign xor_ln302_310_fu_40572_p2 = (xor_ln302_309_fu_40566_p2 ^ 1'd1);

assign xor_ln302_311_fu_40668_p2 = (p_Result_796_fu_40636_p3 ^ p_Result_795_fu_40622_p3);

assign xor_ln302_312_fu_40674_p2 = (xor_ln302_311_fu_40668_p2 ^ 1'd1);

assign xor_ln302_313_fu_40770_p2 = (p_Result_798_fu_40738_p3 ^ p_Result_797_fu_40724_p3);

assign xor_ln302_314_fu_40776_p2 = (xor_ln302_313_fu_40770_p2 ^ 1'd1);

assign xor_ln302_315_fu_40872_p2 = (p_Result_800_fu_40840_p3 ^ p_Result_799_fu_40826_p3);

assign xor_ln302_316_fu_40878_p2 = (xor_ln302_315_fu_40872_p2 ^ 1'd1);

assign xor_ln302_317_fu_40974_p2 = (p_Result_802_fu_40942_p3 ^ p_Result_801_fu_40928_p3);

assign xor_ln302_318_fu_40980_p2 = (xor_ln302_317_fu_40974_p2 ^ 1'd1);

assign xor_ln302_319_fu_41076_p2 = (p_Result_804_fu_41044_p3 ^ p_Result_803_fu_41030_p3);

assign xor_ln302_320_fu_41082_p2 = (xor_ln302_319_fu_41076_p2 ^ 1'd1);

assign xor_ln302_321_fu_41178_p2 = (p_Result_806_fu_41146_p3 ^ p_Result_805_fu_41132_p3);

assign xor_ln302_322_fu_41184_p2 = (xor_ln302_321_fu_41178_p2 ^ 1'd1);

assign xor_ln302_fu_23678_p2 = (p_Result_646_fu_23646_p3 ^ p_Result_645_fu_23632_p3);

assign xor_ln888_160_fu_19104_p2 = (p_Result_406_reg_41370 ^ 1'd1);

assign xor_ln888_162_fu_19229_p2 = (p_Result_409_reg_41401 ^ 1'd1);

assign xor_ln888_164_fu_19354_p2 = (p_Result_412_reg_41432 ^ 1'd1);

assign xor_ln888_166_fu_19479_p2 = (p_Result_415_reg_41463 ^ 1'd1);

assign xor_ln888_168_fu_19604_p2 = (p_Result_418_reg_41494 ^ 1'd1);

assign xor_ln888_170_fu_19729_p2 = (p_Result_421_reg_41525 ^ 1'd1);

assign xor_ln888_172_fu_19854_p2 = (p_Result_424_reg_41556 ^ 1'd1);

assign xor_ln888_174_fu_19979_p2 = (p_Result_427_reg_41587 ^ 1'd1);

assign xor_ln888_176_fu_20126_p2 = (p_Result_430_reg_41623 ^ 1'd1);

assign xor_ln888_178_fu_20275_p2 = (p_Result_433_reg_41652 ^ 1'd1);

assign xor_ln888_180_fu_20424_p2 = (p_Result_436_reg_41681 ^ 1'd1);

assign xor_ln888_182_fu_20573_p2 = (p_Result_439_reg_41710 ^ 1'd1);

assign xor_ln888_184_fu_20722_p2 = (p_Result_442_reg_41739 ^ 1'd1);

assign xor_ln888_186_fu_18203_p2 = (p_Result_445_fu_18149_p3 ^ 1'd1);

assign xor_ln888_188_fu_20888_p2 = (p_Result_448_reg_41783 ^ 1'd1);

assign xor_ln888_190_fu_21037_p2 = (p_Result_451_reg_41812 ^ 1'd1);

assign xor_ln888_192_fu_21186_p2 = (p_Result_454_reg_41841 ^ 1'd1);

assign xor_ln888_194_fu_21331_p2 = (p_Result_457_reg_41870 ^ 1'd1);

assign xor_ln888_196_fu_21476_p2 = (p_Result_460_reg_41899 ^ 1'd1);

assign xor_ln888_198_fu_21605_p2 = (p_Result_463_reg_41928 ^ 1'd1);

assign xor_ln888_200_fu_21730_p2 = (p_Result_466_reg_41957 ^ 1'd1);

assign xor_ln888_202_fu_21875_p2 = (p_Result_469_reg_41986 ^ 1'd1);

assign xor_ln888_204_fu_22004_p2 = (p_Result_472_reg_42015 ^ 1'd1);

assign xor_ln888_206_fu_22133_p2 = (p_Result_475_reg_42044 ^ 1'd1);

assign xor_ln888_208_fu_22262_p2 = (p_Result_478_reg_42073 ^ 1'd1);

assign xor_ln888_210_fu_22391_p2 = (p_Result_481_reg_42102 ^ 1'd1);

assign xor_ln888_212_fu_25554_p2 = (p_Result_484_reg_42258 ^ 1'd1);

assign xor_ln888_214_fu_25679_p2 = (p_Result_487_reg_42289 ^ 1'd1);

assign xor_ln888_216_fu_25804_p2 = (p_Result_490_reg_42320 ^ 1'd1);

assign xor_ln888_218_fu_25929_p2 = (p_Result_493_reg_42351 ^ 1'd1);

assign xor_ln888_220_fu_26054_p2 = (p_Result_496_reg_42382 ^ 1'd1);

assign xor_ln888_222_fu_26179_p2 = (p_Result_499_reg_42413 ^ 1'd1);

assign xor_ln888_224_fu_22985_p2 = (p_Result_502_fu_22940_p3 ^ 1'd1);

assign xor_ln888_226_fu_26321_p2 = (p_Result_505_reg_42459 ^ 1'd1);

assign xor_ln888_228_fu_26446_p2 = (p_Result_508_reg_42490 ^ 1'd1);

assign xor_ln888_230_fu_26589_p2 = (p_Result_511_reg_42526 ^ 1'd1);

assign xor_ln888_232_fu_26738_p2 = (p_Result_514_reg_42555 ^ 1'd1);

assign xor_ln888_234_fu_26887_p2 = (p_Result_517_reg_42584 ^ 1'd1);

assign xor_ln888_236_fu_27036_p2 = (p_Result_520_reg_42613 ^ 1'd1);

assign xor_ln888_238_fu_27185_p2 = (p_Result_523_reg_42642 ^ 1'd1);

assign xor_ln888_240_fu_27334_p2 = (p_Result_526_reg_42671 ^ 1'd1);

assign xor_ln888_242_fu_27483_p2 = (p_Result_529_reg_42700 ^ 1'd1);

assign xor_ln888_244_fu_27632_p2 = (p_Result_532_reg_42729 ^ 1'd1);

assign xor_ln888_246_fu_27781_p2 = (p_Result_535_reg_42758 ^ 1'd1);

assign xor_ln888_248_fu_28013_p2 = (p_Result_538_fu_27968_p3 ^ 1'd1);

assign xor_ln888_250_fu_31352_p2 = (p_Result_541_reg_42851 ^ 1'd1);

assign xor_ln888_252_fu_31477_p2 = (p_Result_544_reg_42882 ^ 1'd1);

assign xor_ln888_254_fu_31602_p2 = (p_Result_547_reg_42913 ^ 1'd1);

assign xor_ln888_256_fu_31727_p2 = (p_Result_550_reg_42944 ^ 1'd1);

assign xor_ln888_258_fu_31852_p2 = (p_Result_553_reg_42975 ^ 1'd1);

assign xor_ln888_260_fu_31977_p2 = (p_Result_556_reg_43006 ^ 1'd1);

assign xor_ln888_262_fu_32102_p2 = (p_Result_559_reg_43037 ^ 1'd1);

assign xor_ln888_264_fu_32227_p2 = (p_Result_562_reg_43068 ^ 1'd1);

assign xor_ln888_266_fu_32374_p2 = (p_Result_565_reg_43104 ^ 1'd1);

assign xor_ln888_268_fu_32523_p2 = (p_Result_568_reg_43133 ^ 1'd1);

assign xor_ln888_270_fu_32672_p2 = (p_Result_571_reg_43162 ^ 1'd1);

assign xor_ln888_272_fu_32821_p2 = (p_Result_574_reg_43191 ^ 1'd1);

assign xor_ln888_274_fu_32970_p2 = (p_Result_577_reg_43220 ^ 1'd1);

assign xor_ln888_276_fu_33119_p2 = (p_Result_580_reg_43249 ^ 1'd1);

assign xor_ln888_278_fu_33268_p2 = (p_Result_583_reg_43278 ^ 1'd1);

assign xor_ln888_280_fu_33417_p2 = (p_Result_586_reg_43307 ^ 1'd1);

assign xor_ln888_282_fu_29080_p2 = (p_Result_589_fu_29035_p3 ^ 1'd1);

assign xor_ln888_284_fu_37086_p2 = (p_Result_592_reg_43526 ^ 1'd1);

assign xor_ln888_286_fu_37210_p2 = (p_Result_595_reg_43557 ^ 1'd1);

assign xor_ln888_288_fu_37335_p2 = (p_Result_598_reg_43588 ^ 1'd1);

assign xor_ln888_290_fu_37460_p2 = (p_Result_601_reg_43619 ^ 1'd1);

assign xor_ln888_292_fu_37585_p2 = (p_Result_604_reg_43650 ^ 1'd1);

assign xor_ln888_294_fu_37710_p2 = (p_Result_607_reg_43681 ^ 1'd1);

assign xor_ln888_296_fu_37835_p2 = (p_Result_610_reg_43712 ^ 1'd1);

assign xor_ln888_298_fu_37960_p2 = (p_Result_613_reg_43743 ^ 1'd1);

assign xor_ln888_300_fu_38085_p2 = (p_Result_616_reg_43774 ^ 1'd1);

assign xor_ln888_302_fu_38228_p2 = (p_Result_619_reg_43810 ^ 1'd1);

assign xor_ln888_304_fu_38377_p2 = (p_Result_622_reg_43839 ^ 1'd1);

assign xor_ln888_306_fu_38526_p2 = (p_Result_625_reg_43868 ^ 1'd1);

assign xor_ln888_308_fu_38675_p2 = (p_Result_628_reg_43897 ^ 1'd1);

assign xor_ln888_310_fu_38824_p2 = (p_Result_631_reg_43926 ^ 1'd1);

assign xor_ln888_312_fu_38973_p2 = (p_Result_634_reg_43955 ^ 1'd1);

assign xor_ln888_314_fu_39122_p2 = (p_Result_637_reg_43984 ^ 1'd1);

assign xor_ln888_316_fu_34572_p2 = (p_Result_640_fu_34518_p3 ^ 1'd1);

assign xor_ln888_318_fu_39288_p2 = (p_Result_643_reg_44028 ^ 1'd1);

assign xor_ln888_fu_18979_p2 = (p_Result_403_reg_41339 ^ 1'd1);

assign xor_ln890_100_fu_21899_p2 = (tmp_774_fu_21891_p3 ^ 1'd1);

assign xor_ln890_101_fu_22028_p2 = (tmp_780_fu_22020_p3 ^ 1'd1);

assign xor_ln890_102_fu_22157_p2 = (tmp_786_fu_22149_p3 ^ 1'd1);

assign xor_ln890_103_fu_22286_p2 = (tmp_792_fu_22278_p3 ^ 1'd1);

assign xor_ln890_104_fu_22415_p2 = (tmp_798_fu_22407_p3 ^ 1'd1);

assign xor_ln890_105_fu_25577_p2 = (tmp_804_fu_25569_p3 ^ 1'd1);

assign xor_ln890_106_fu_25702_p2 = (tmp_810_fu_25694_p3 ^ 1'd1);

assign xor_ln890_107_fu_25827_p2 = (tmp_816_fu_25819_p3 ^ 1'd1);

assign xor_ln890_108_fu_25952_p2 = (tmp_822_fu_25944_p3 ^ 1'd1);

assign xor_ln890_109_fu_26077_p2 = (tmp_828_fu_26069_p3 ^ 1'd1);

assign xor_ln890_110_fu_26202_p2 = (tmp_834_fu_26194_p3 ^ 1'd1);

assign xor_ln890_111_fu_23011_p2 = (tmp_840_fu_23003_p3 ^ 1'd1);

assign xor_ln890_112_fu_26344_p2 = (tmp_846_fu_26336_p3 ^ 1'd1);

assign xor_ln890_113_fu_26469_p2 = (tmp_852_fu_26461_p3 ^ 1'd1);

assign xor_ln890_114_fu_26613_p2 = (tmp_858_fu_26605_p3 ^ 1'd1);

assign xor_ln890_115_fu_26762_p2 = (tmp_864_fu_26754_p3 ^ 1'd1);

assign xor_ln890_116_fu_26911_p2 = (tmp_870_fu_26903_p3 ^ 1'd1);

assign xor_ln890_117_fu_27060_p2 = (tmp_876_fu_27052_p3 ^ 1'd1);

assign xor_ln890_118_fu_27209_p2 = (tmp_882_fu_27201_p3 ^ 1'd1);

assign xor_ln890_119_fu_27358_p2 = (tmp_888_fu_27350_p3 ^ 1'd1);

assign xor_ln890_120_fu_27507_p2 = (tmp_894_fu_27499_p3 ^ 1'd1);

assign xor_ln890_121_fu_27656_p2 = (tmp_900_fu_27648_p3 ^ 1'd1);

assign xor_ln890_122_fu_27805_p2 = (tmp_906_fu_27797_p3 ^ 1'd1);

assign xor_ln890_123_fu_28039_p2 = (tmp_912_fu_28031_p3 ^ 1'd1);

assign xor_ln890_124_fu_31375_p2 = (tmp_918_fu_31367_p3 ^ 1'd1);

assign xor_ln890_125_fu_31500_p2 = (tmp_924_fu_31492_p3 ^ 1'd1);

assign xor_ln890_126_fu_31625_p2 = (tmp_930_fu_31617_p3 ^ 1'd1);

assign xor_ln890_127_fu_31750_p2 = (tmp_936_fu_31742_p3 ^ 1'd1);

assign xor_ln890_128_fu_31875_p2 = (tmp_942_fu_31867_p3 ^ 1'd1);

assign xor_ln890_129_fu_32000_p2 = (tmp_948_fu_31992_p3 ^ 1'd1);

assign xor_ln890_130_fu_32125_p2 = (tmp_954_fu_32117_p3 ^ 1'd1);

assign xor_ln890_131_fu_32250_p2 = (tmp_960_fu_32242_p3 ^ 1'd1);

assign xor_ln890_132_fu_32398_p2 = (tmp_966_fu_32390_p3 ^ 1'd1);

assign xor_ln890_133_fu_32547_p2 = (tmp_972_fu_32539_p3 ^ 1'd1);

assign xor_ln890_134_fu_32696_p2 = (tmp_978_fu_32688_p3 ^ 1'd1);

assign xor_ln890_135_fu_32845_p2 = (tmp_984_fu_32837_p3 ^ 1'd1);

assign xor_ln890_136_fu_32994_p2 = (tmp_990_fu_32986_p3 ^ 1'd1);

assign xor_ln890_137_fu_33143_p2 = (tmp_996_fu_33135_p3 ^ 1'd1);

assign xor_ln890_138_fu_33292_p2 = (tmp_1002_fu_33284_p3 ^ 1'd1);

assign xor_ln890_139_fu_33441_p2 = (tmp_1008_fu_33433_p3 ^ 1'd1);

assign xor_ln890_140_fu_29106_p2 = (tmp_1014_fu_29098_p3 ^ 1'd1);

assign xor_ln890_141_fu_37109_p2 = (tmp_1020_fu_37101_p3 ^ 1'd1);

assign xor_ln890_142_fu_37233_p2 = (tmp_1026_fu_37225_p3 ^ 1'd1);

assign xor_ln890_143_fu_37358_p2 = (tmp_1032_fu_37350_p3 ^ 1'd1);

assign xor_ln890_144_fu_37483_p2 = (tmp_1038_fu_37475_p3 ^ 1'd1);

assign xor_ln890_145_fu_37608_p2 = (tmp_1044_fu_37600_p3 ^ 1'd1);

assign xor_ln890_146_fu_37733_p2 = (tmp_1050_fu_37725_p3 ^ 1'd1);

assign xor_ln890_147_fu_37858_p2 = (tmp_1056_fu_37850_p3 ^ 1'd1);

assign xor_ln890_148_fu_37983_p2 = (tmp_1062_fu_37975_p3 ^ 1'd1);

assign xor_ln890_149_fu_38108_p2 = (tmp_1068_fu_38100_p3 ^ 1'd1);

assign xor_ln890_150_fu_38252_p2 = (tmp_1074_fu_38244_p3 ^ 1'd1);

assign xor_ln890_151_fu_38401_p2 = (tmp_1080_fu_38393_p3 ^ 1'd1);

assign xor_ln890_152_fu_38550_p2 = (tmp_1086_fu_38542_p3 ^ 1'd1);

assign xor_ln890_153_fu_38699_p2 = (tmp_1092_fu_38691_p3 ^ 1'd1);

assign xor_ln890_154_fu_38848_p2 = (tmp_1098_fu_38840_p3 ^ 1'd1);

assign xor_ln890_155_fu_38997_p2 = (tmp_1104_fu_38989_p3 ^ 1'd1);

assign xor_ln890_156_fu_39146_p2 = (tmp_1110_fu_39138_p3 ^ 1'd1);

assign xor_ln890_157_fu_34598_p2 = (tmp_1116_fu_34590_p3 ^ 1'd1);

assign xor_ln890_158_fu_39312_p2 = (tmp_1122_fu_39304_p3 ^ 1'd1);

assign xor_ln890_79_fu_19127_p2 = (tmp_648_fu_19119_p3 ^ 1'd1);

assign xor_ln890_80_fu_19252_p2 = (tmp_654_fu_19244_p3 ^ 1'd1);

assign xor_ln890_81_fu_19377_p2 = (tmp_660_fu_19369_p3 ^ 1'd1);

assign xor_ln890_82_fu_19502_p2 = (tmp_666_fu_19494_p3 ^ 1'd1);

assign xor_ln890_83_fu_19627_p2 = (tmp_672_fu_19619_p3 ^ 1'd1);

assign xor_ln890_84_fu_19752_p2 = (tmp_678_fu_19744_p3 ^ 1'd1);

assign xor_ln890_85_fu_19877_p2 = (tmp_684_fu_19869_p3 ^ 1'd1);

assign xor_ln890_86_fu_20002_p2 = (tmp_690_fu_19994_p3 ^ 1'd1);

assign xor_ln890_87_fu_20150_p2 = (tmp_696_fu_20142_p3 ^ 1'd1);

assign xor_ln890_88_fu_20299_p2 = (tmp_702_fu_20291_p3 ^ 1'd1);

assign xor_ln890_89_fu_20448_p2 = (tmp_708_fu_20440_p3 ^ 1'd1);

assign xor_ln890_90_fu_20597_p2 = (tmp_714_fu_20589_p3 ^ 1'd1);

assign xor_ln890_91_fu_20746_p2 = (tmp_720_fu_20738_p3 ^ 1'd1);

assign xor_ln890_92_fu_18229_p2 = (tmp_726_fu_18221_p3 ^ 1'd1);

assign xor_ln890_93_fu_20912_p2 = (tmp_732_fu_20904_p3 ^ 1'd1);

assign xor_ln890_94_fu_21061_p2 = (tmp_738_fu_21053_p3 ^ 1'd1);

assign xor_ln890_95_fu_21210_p2 = (tmp_744_fu_21202_p3 ^ 1'd1);

assign xor_ln890_96_fu_21355_p2 = (tmp_750_fu_21347_p3 ^ 1'd1);

assign xor_ln890_97_fu_21500_p2 = (tmp_756_fu_21492_p3 ^ 1'd1);

assign xor_ln890_98_fu_21629_p2 = (tmp_762_fu_21621_p3 ^ 1'd1);

assign xor_ln890_99_fu_21754_p2 = (tmp_768_fu_21746_p3 ^ 1'd1);

assign xor_ln890_fu_19002_p2 = (tmp_642_fu_18994_p3 ^ 1'd1);

assign xor_ln895_243_fu_19035_p2 = (p_Result_s_reg_41333 ^ 1'd1);

assign xor_ln895_244_fu_19149_p2 = (deleted_zeros_78_fu_19114_p2 ^ 1'd1);

assign xor_ln895_245_fu_19160_p2 = (p_Result_405_reg_41364 ^ 1'd1);

assign xor_ln895_246_fu_19274_p2 = (deleted_zeros_79_fu_19239_p2 ^ 1'd1);

assign xor_ln895_247_fu_19285_p2 = (p_Result_408_reg_41395 ^ 1'd1);

assign xor_ln895_248_fu_19399_p2 = (deleted_zeros_80_fu_19364_p2 ^ 1'd1);

assign xor_ln895_249_fu_19410_p2 = (p_Result_411_reg_41426 ^ 1'd1);

assign xor_ln895_250_fu_19524_p2 = (deleted_zeros_81_fu_19489_p2 ^ 1'd1);

assign xor_ln895_251_fu_19535_p2 = (p_Result_414_reg_41457 ^ 1'd1);

assign xor_ln895_252_fu_19649_p2 = (deleted_zeros_82_fu_19614_p2 ^ 1'd1);

assign xor_ln895_253_fu_19660_p2 = (p_Result_417_reg_41488 ^ 1'd1);

assign xor_ln895_254_fu_19774_p2 = (deleted_zeros_83_fu_19739_p2 ^ 1'd1);

assign xor_ln895_255_fu_19785_p2 = (p_Result_420_reg_41519 ^ 1'd1);

assign xor_ln895_256_fu_19899_p2 = (deleted_zeros_84_fu_19864_p2 ^ 1'd1);

assign xor_ln895_257_fu_19910_p2 = (p_Result_423_reg_41550 ^ 1'd1);

assign xor_ln895_258_fu_20024_p2 = (deleted_zeros_85_fu_19989_p2 ^ 1'd1);

assign xor_ln895_259_fu_20035_p2 = (p_Result_426_reg_41581 ^ 1'd1);

assign xor_ln895_260_fu_20172_p2 = (deleted_zeros_86_fu_20137_p2 ^ 1'd1);

assign xor_ln895_261_fu_20184_p2 = (p_Result_429_reg_41612 ^ 1'd1);

assign xor_ln895_262_fu_20321_p2 = (deleted_zeros_87_fu_20286_p2 ^ 1'd1);

assign xor_ln895_263_fu_20333_p2 = (p_Result_432_reg_41641 ^ 1'd1);

assign xor_ln895_264_fu_20470_p2 = (deleted_zeros_88_fu_20435_p2 ^ 1'd1);

assign xor_ln895_265_fu_20482_p2 = (p_Result_435_reg_41670 ^ 1'd1);

assign xor_ln895_266_fu_20619_p2 = (deleted_zeros_89_fu_20584_p2 ^ 1'd1);

assign xor_ln895_267_fu_20631_p2 = (p_Result_438_reg_41699 ^ 1'd1);

assign xor_ln895_268_fu_20768_p2 = (deleted_zeros_90_fu_20733_p2 ^ 1'd1);

assign xor_ln895_269_fu_20780_p2 = (p_Result_441_reg_41728 ^ 1'd1);

assign xor_ln895_270_fu_18253_p2 = (deleted_zeros_91_fu_18215_p2 ^ 1'd1);

assign xor_ln895_271_fu_18265_p2 = (p_Result_444_fu_18127_p3 ^ 1'd1);

assign xor_ln895_272_fu_20934_p2 = (deleted_zeros_92_fu_20899_p2 ^ 1'd1);

assign xor_ln895_273_fu_20946_p2 = (p_Result_447_reg_41772 ^ 1'd1);

assign xor_ln895_274_fu_21083_p2 = (deleted_zeros_93_fu_21048_p2 ^ 1'd1);

assign xor_ln895_275_fu_21095_p2 = (p_Result_450_reg_41801 ^ 1'd1);

assign xor_ln895_276_fu_21232_p2 = (deleted_zeros_94_fu_21197_p2 ^ 1'd1);

assign xor_ln895_277_fu_21244_p2 = (p_Result_453_reg_41830 ^ 1'd1);

assign xor_ln895_278_fu_21377_p2 = (deleted_zeros_95_fu_21342_p2 ^ 1'd1);

assign xor_ln895_279_fu_21389_p2 = (p_Result_456_reg_41859 ^ 1'd1);

assign xor_ln895_280_fu_21522_p2 = (deleted_zeros_96_fu_21487_p2 ^ 1'd1);

assign xor_ln895_281_fu_21534_p2 = (p_Result_459_reg_41888 ^ 1'd1);

assign xor_ln895_282_fu_21651_p2 = (deleted_zeros_97_fu_21616_p2 ^ 1'd1);

assign xor_ln895_283_fu_21663_p2 = (p_Result_462_reg_41917 ^ 1'd1);

assign xor_ln895_284_fu_21776_p2 = (deleted_zeros_98_fu_21741_p2 ^ 1'd1);

assign xor_ln895_285_fu_21788_p2 = (p_Result_465_reg_41946 ^ 1'd1);

assign xor_ln895_286_fu_21921_p2 = (deleted_zeros_99_fu_21886_p2 ^ 1'd1);

assign xor_ln895_287_fu_21933_p2 = (p_Result_468_reg_41975 ^ 1'd1);

assign xor_ln895_288_fu_22050_p2 = (deleted_zeros_100_fu_22015_p2 ^ 1'd1);

assign xor_ln895_289_fu_22062_p2 = (p_Result_471_reg_42004 ^ 1'd1);

assign xor_ln895_290_fu_22179_p2 = (deleted_zeros_101_fu_22144_p2 ^ 1'd1);

assign xor_ln895_291_fu_22191_p2 = (p_Result_474_reg_42033 ^ 1'd1);

assign xor_ln895_292_fu_22308_p2 = (deleted_zeros_102_fu_22273_p2 ^ 1'd1);

assign xor_ln895_293_fu_22320_p2 = (p_Result_477_reg_42062 ^ 1'd1);

assign xor_ln895_294_fu_22437_p2 = (deleted_zeros_103_fu_22402_p2 ^ 1'd1);

assign xor_ln895_295_fu_22449_p2 = (p_Result_480_reg_42091 ^ 1'd1);

assign xor_ln895_296_fu_25599_p2 = (deleted_zeros_104_fu_25564_p2 ^ 1'd1);

assign xor_ln895_297_fu_25610_p2 = (p_Result_483_reg_42252 ^ 1'd1);

assign xor_ln895_298_fu_25724_p2 = (deleted_zeros_105_fu_25689_p2 ^ 1'd1);

assign xor_ln895_299_fu_25735_p2 = (p_Result_486_reg_42283 ^ 1'd1);

assign xor_ln895_300_fu_25849_p2 = (deleted_zeros_106_fu_25814_p2 ^ 1'd1);

assign xor_ln895_301_fu_25860_p2 = (p_Result_489_reg_42314 ^ 1'd1);

assign xor_ln895_302_fu_25974_p2 = (deleted_zeros_107_fu_25939_p2 ^ 1'd1);

assign xor_ln895_303_fu_25985_p2 = (p_Result_492_reg_42345 ^ 1'd1);

assign xor_ln895_304_fu_26099_p2 = (deleted_zeros_108_fu_26064_p2 ^ 1'd1);

assign xor_ln895_305_fu_26110_p2 = (p_Result_495_reg_42376 ^ 1'd1);

assign xor_ln895_306_fu_26224_p2 = (deleted_zeros_109_fu_26189_p2 ^ 1'd1);

assign xor_ln895_307_fu_26235_p2 = (p_Result_498_reg_42407 ^ 1'd1);

assign xor_ln895_308_fu_23035_p2 = (deleted_zeros_110_fu_22997_p2 ^ 1'd1);

assign xor_ln895_309_fu_23047_p2 = (p_Result_501_fu_22918_p3 ^ 1'd1);

assign xor_ln895_310_fu_26366_p2 = (deleted_zeros_111_fu_26331_p2 ^ 1'd1);

assign xor_ln895_311_fu_26377_p2 = (p_Result_504_reg_42453 ^ 1'd1);

assign xor_ln895_312_fu_26491_p2 = (deleted_zeros_112_fu_26456_p2 ^ 1'd1);

assign xor_ln895_313_fu_26502_p2 = (p_Result_507_reg_42484 ^ 1'd1);

assign xor_ln895_314_fu_26635_p2 = (deleted_zeros_113_fu_26600_p2 ^ 1'd1);

assign xor_ln895_315_fu_26647_p2 = (p_Result_510_reg_42515 ^ 1'd1);

assign xor_ln895_316_fu_26784_p2 = (deleted_zeros_114_fu_26749_p2 ^ 1'd1);

assign xor_ln895_317_fu_26796_p2 = (p_Result_513_reg_42544 ^ 1'd1);

assign xor_ln895_318_fu_26933_p2 = (deleted_zeros_115_fu_26898_p2 ^ 1'd1);

assign xor_ln895_319_fu_26945_p2 = (p_Result_516_reg_42573 ^ 1'd1);

assign xor_ln895_320_fu_27082_p2 = (deleted_zeros_116_fu_27047_p2 ^ 1'd1);

assign xor_ln895_321_fu_27094_p2 = (p_Result_519_reg_42602 ^ 1'd1);

assign xor_ln895_322_fu_27231_p2 = (deleted_zeros_117_fu_27196_p2 ^ 1'd1);

assign xor_ln895_323_fu_27243_p2 = (p_Result_522_reg_42631 ^ 1'd1);

assign xor_ln895_324_fu_27380_p2 = (deleted_zeros_118_fu_27345_p2 ^ 1'd1);

assign xor_ln895_325_fu_27392_p2 = (p_Result_525_reg_42660 ^ 1'd1);

assign xor_ln895_326_fu_27529_p2 = (deleted_zeros_119_fu_27494_p2 ^ 1'd1);

assign xor_ln895_327_fu_27541_p2 = (p_Result_528_reg_42689 ^ 1'd1);

assign xor_ln895_328_fu_27678_p2 = (deleted_zeros_120_fu_27643_p2 ^ 1'd1);

assign xor_ln895_329_fu_27690_p2 = (p_Result_531_reg_42718 ^ 1'd1);

assign xor_ln895_330_fu_27827_p2 = (deleted_zeros_121_fu_27792_p2 ^ 1'd1);

assign xor_ln895_331_fu_27839_p2 = (p_Result_534_reg_42747 ^ 1'd1);

assign xor_ln895_332_fu_28063_p2 = (deleted_zeros_122_fu_28025_p2 ^ 1'd1);

assign xor_ln895_333_fu_28075_p2 = (p_Result_537_fu_27946_p3 ^ 1'd1);

assign xor_ln895_334_fu_31397_p2 = (deleted_zeros_123_fu_31362_p2 ^ 1'd1);

assign xor_ln895_335_fu_31408_p2 = (p_Result_540_reg_42845 ^ 1'd1);

assign xor_ln895_336_fu_31522_p2 = (deleted_zeros_124_fu_31487_p2 ^ 1'd1);

assign xor_ln895_337_fu_31533_p2 = (p_Result_543_reg_42876 ^ 1'd1);

assign xor_ln895_338_fu_31647_p2 = (deleted_zeros_125_fu_31612_p2 ^ 1'd1);

assign xor_ln895_339_fu_31658_p2 = (p_Result_546_reg_42907 ^ 1'd1);

assign xor_ln895_340_fu_31772_p2 = (deleted_zeros_126_fu_31737_p2 ^ 1'd1);

assign xor_ln895_341_fu_31783_p2 = (p_Result_549_reg_42938 ^ 1'd1);

assign xor_ln895_342_fu_31897_p2 = (deleted_zeros_127_fu_31862_p2 ^ 1'd1);

assign xor_ln895_343_fu_31908_p2 = (p_Result_552_reg_42969 ^ 1'd1);

assign xor_ln895_344_fu_32022_p2 = (deleted_zeros_128_fu_31987_p2 ^ 1'd1);

assign xor_ln895_345_fu_32033_p2 = (p_Result_555_reg_43000 ^ 1'd1);

assign xor_ln895_346_fu_32147_p2 = (deleted_zeros_129_fu_32112_p2 ^ 1'd1);

assign xor_ln895_347_fu_32158_p2 = (p_Result_558_reg_43031 ^ 1'd1);

assign xor_ln895_348_fu_32272_p2 = (deleted_zeros_130_fu_32237_p2 ^ 1'd1);

assign xor_ln895_349_fu_32283_p2 = (p_Result_561_reg_43062 ^ 1'd1);

assign xor_ln895_350_fu_32420_p2 = (deleted_zeros_131_fu_32385_p2 ^ 1'd1);

assign xor_ln895_351_fu_32432_p2 = (p_Result_564_reg_43093 ^ 1'd1);

assign xor_ln895_352_fu_32569_p2 = (deleted_zeros_132_fu_32534_p2 ^ 1'd1);

assign xor_ln895_353_fu_32581_p2 = (p_Result_567_reg_43122 ^ 1'd1);

assign xor_ln895_354_fu_32718_p2 = (deleted_zeros_133_fu_32683_p2 ^ 1'd1);

assign xor_ln895_355_fu_32730_p2 = (p_Result_570_reg_43151 ^ 1'd1);

assign xor_ln895_356_fu_32867_p2 = (deleted_zeros_134_fu_32832_p2 ^ 1'd1);

assign xor_ln895_357_fu_32879_p2 = (p_Result_573_reg_43180 ^ 1'd1);

assign xor_ln895_358_fu_33016_p2 = (deleted_zeros_135_fu_32981_p2 ^ 1'd1);

assign xor_ln895_359_fu_33028_p2 = (p_Result_576_reg_43209 ^ 1'd1);

assign xor_ln895_360_fu_33165_p2 = (deleted_zeros_136_fu_33130_p2 ^ 1'd1);

assign xor_ln895_361_fu_33177_p2 = (p_Result_579_reg_43238 ^ 1'd1);

assign xor_ln895_362_fu_33314_p2 = (deleted_zeros_137_fu_33279_p2 ^ 1'd1);

assign xor_ln895_363_fu_33326_p2 = (p_Result_582_reg_43267 ^ 1'd1);

assign xor_ln895_364_fu_33463_p2 = (deleted_zeros_138_fu_33428_p2 ^ 1'd1);

assign xor_ln895_365_fu_33475_p2 = (p_Result_585_reg_43296 ^ 1'd1);

assign xor_ln895_366_fu_29130_p2 = (deleted_zeros_139_fu_29092_p2 ^ 1'd1);

assign xor_ln895_367_fu_29142_p2 = (p_Result_588_fu_29013_p3 ^ 1'd1);

assign xor_ln895_368_fu_37131_p2 = (deleted_zeros_140_fu_37096_p2 ^ 1'd1);

assign xor_ln895_369_fu_37142_p2 = (p_Result_591_reg_43520 ^ 1'd1);

assign xor_ln895_370_fu_37255_p2 = (deleted_zeros_141_fu_37220_p2 ^ 1'd1);

assign xor_ln895_371_fu_37266_p2 = (p_Result_594_reg_43551 ^ 1'd1);

assign xor_ln895_372_fu_37380_p2 = (deleted_zeros_142_fu_37345_p2 ^ 1'd1);

assign xor_ln895_373_fu_37391_p2 = (p_Result_597_reg_43582 ^ 1'd1);

assign xor_ln895_374_fu_37505_p2 = (deleted_zeros_143_fu_37470_p2 ^ 1'd1);

assign xor_ln895_375_fu_37516_p2 = (p_Result_600_reg_43613 ^ 1'd1);

assign xor_ln895_376_fu_37630_p2 = (deleted_zeros_144_fu_37595_p2 ^ 1'd1);

assign xor_ln895_377_fu_37641_p2 = (p_Result_603_reg_43644 ^ 1'd1);

assign xor_ln895_378_fu_37755_p2 = (deleted_zeros_145_fu_37720_p2 ^ 1'd1);

assign xor_ln895_379_fu_37766_p2 = (p_Result_606_reg_43675 ^ 1'd1);

assign xor_ln895_380_fu_37880_p2 = (deleted_zeros_146_fu_37845_p2 ^ 1'd1);

assign xor_ln895_381_fu_37891_p2 = (p_Result_609_reg_43706 ^ 1'd1);

assign xor_ln895_382_fu_38005_p2 = (deleted_zeros_147_fu_37970_p2 ^ 1'd1);

assign xor_ln895_383_fu_38016_p2 = (p_Result_612_reg_43737 ^ 1'd1);

assign xor_ln895_384_fu_38130_p2 = (deleted_zeros_148_fu_38095_p2 ^ 1'd1);

assign xor_ln895_385_fu_38141_p2 = (p_Result_615_reg_43768 ^ 1'd1);

assign xor_ln895_386_fu_38274_p2 = (deleted_zeros_149_fu_38239_p2 ^ 1'd1);

assign xor_ln895_387_fu_38286_p2 = (p_Result_618_reg_43799 ^ 1'd1);

assign xor_ln895_388_fu_38423_p2 = (deleted_zeros_150_fu_38388_p2 ^ 1'd1);

assign xor_ln895_389_fu_38435_p2 = (p_Result_621_reg_43828 ^ 1'd1);

assign xor_ln895_390_fu_38572_p2 = (deleted_zeros_151_fu_38537_p2 ^ 1'd1);

assign xor_ln895_391_fu_38584_p2 = (p_Result_624_reg_43857 ^ 1'd1);

assign xor_ln895_392_fu_38721_p2 = (deleted_zeros_152_fu_38686_p2 ^ 1'd1);

assign xor_ln895_393_fu_38733_p2 = (p_Result_627_reg_43886 ^ 1'd1);

assign xor_ln895_394_fu_38870_p2 = (deleted_zeros_153_fu_38835_p2 ^ 1'd1);

assign xor_ln895_395_fu_38882_p2 = (p_Result_630_reg_43915 ^ 1'd1);

assign xor_ln895_396_fu_39019_p2 = (deleted_zeros_154_fu_38984_p2 ^ 1'd1);

assign xor_ln895_397_fu_39031_p2 = (p_Result_633_reg_43944 ^ 1'd1);

assign xor_ln895_398_fu_39168_p2 = (deleted_zeros_155_fu_39133_p2 ^ 1'd1);

assign xor_ln895_399_fu_39180_p2 = (p_Result_636_reg_43973 ^ 1'd1);

assign xor_ln895_400_fu_34622_p2 = (deleted_zeros_156_fu_34584_p2 ^ 1'd1);

assign xor_ln895_401_fu_34634_p2 = (p_Result_639_fu_34496_p3 ^ 1'd1);

assign xor_ln895_402_fu_39334_p2 = (deleted_zeros_157_fu_39299_p2 ^ 1'd1);

assign xor_ln895_403_fu_39346_p2 = (p_Result_642_reg_44017 ^ 1'd1);

assign xor_ln895_404_fu_23654_p2 = (p_Result_645_fu_23632_p3 ^ 1'd1);

assign xor_ln895_405_fu_23752_p2 = (p_Result_647_fu_23730_p3 ^ 1'd1);

assign xor_ln895_406_fu_23850_p2 = (p_Result_649_fu_23828_p3 ^ 1'd1);

assign xor_ln895_407_fu_23948_p2 = (p_Result_651_fu_23926_p3 ^ 1'd1);

assign xor_ln895_408_fu_24046_p2 = (p_Result_653_fu_24024_p3 ^ 1'd1);

assign xor_ln895_409_fu_24144_p2 = (p_Result_655_fu_24122_p3 ^ 1'd1);

assign xor_ln895_410_fu_24242_p2 = (p_Result_657_fu_24220_p3 ^ 1'd1);

assign xor_ln895_411_fu_24340_p2 = (p_Result_659_fu_24318_p3 ^ 1'd1);

assign xor_ln895_412_fu_24438_p2 = (p_Result_661_fu_24416_p3 ^ 1'd1);

assign xor_ln895_413_fu_24540_p2 = (p_Result_663_fu_24518_p3 ^ 1'd1);

assign xor_ln895_414_fu_24642_p2 = (p_Result_665_fu_24620_p3 ^ 1'd1);

assign xor_ln895_415_fu_24744_p2 = (p_Result_667_fu_24722_p3 ^ 1'd1);

assign xor_ln895_416_fu_24846_p2 = (p_Result_669_fu_24824_p3 ^ 1'd1);

assign xor_ln895_417_fu_24948_p2 = (p_Result_671_fu_24926_p3 ^ 1'd1);

assign xor_ln895_418_fu_25050_p2 = (p_Result_673_fu_25028_p3 ^ 1'd1);

assign xor_ln895_419_fu_25152_p2 = (p_Result_675_fu_25130_p3 ^ 1'd1);

assign xor_ln895_420_fu_25254_p2 = (p_Result_677_fu_25232_p3 ^ 1'd1);

assign xor_ln895_421_fu_25356_p2 = (p_Result_679_fu_25334_p3 ^ 1'd1);

assign xor_ln895_422_fu_29216_p2 = (p_Result_681_fu_29196_p3 ^ 1'd1);

assign xor_ln895_423_fu_29316_p2 = (p_Result_683_fu_29295_p3 ^ 1'd1);

assign xor_ln895_424_fu_29416_p2 = (p_Result_685_fu_29395_p3 ^ 1'd1);

assign xor_ln895_425_fu_29514_p2 = (p_Result_687_fu_29494_p3 ^ 1'd1);

assign xor_ln895_426_fu_29614_p2 = (p_Result_689_fu_29593_p3 ^ 1'd1);

assign xor_ln895_427_fu_29714_p2 = (p_Result_691_fu_29693_p3 ^ 1'd1);

assign xor_ln895_428_fu_29814_p2 = (p_Result_693_fu_29793_p3 ^ 1'd1);

assign xor_ln895_429_fu_29914_p2 = (p_Result_695_fu_29893_p3 ^ 1'd1);

assign xor_ln895_430_fu_30014_p2 = (p_Result_697_fu_29993_p3 ^ 1'd1);

assign xor_ln895_431_fu_30116_p2 = (p_Result_699_fu_30094_p3 ^ 1'd1);

assign xor_ln895_432_fu_30218_p2 = (p_Result_701_fu_30196_p3 ^ 1'd1);

assign xor_ln895_433_fu_30320_p2 = (p_Result_703_fu_30298_p3 ^ 1'd1);

assign xor_ln895_434_fu_30422_p2 = (p_Result_705_fu_30400_p3 ^ 1'd1);

assign xor_ln895_435_fu_30524_p2 = (p_Result_707_fu_30502_p3 ^ 1'd1);

assign xor_ln895_436_fu_30626_p2 = (p_Result_709_fu_30604_p3 ^ 1'd1);

assign xor_ln895_437_fu_30728_p2 = (p_Result_711_fu_30706_p3 ^ 1'd1);

assign xor_ln895_438_fu_30830_p2 = (p_Result_713_fu_30808_p3 ^ 1'd1);

assign xor_ln895_439_fu_30932_p2 = (p_Result_715_fu_30910_p3 ^ 1'd1);

assign xor_ln895_440_fu_34718_p2 = (p_Result_717_reg_43340 ^ 1'd1);

assign xor_ln895_441_fu_34776_p2 = (p_Result_719_reg_43360 ^ 1'd1);

assign xor_ln895_442_fu_34834_p2 = (p_Result_721_reg_43380 ^ 1'd1);

assign xor_ln895_443_fu_34892_p2 = (p_Result_723_reg_43400 ^ 1'd1);

assign xor_ln895_444_fu_34950_p2 = (p_Result_725_reg_43420 ^ 1'd1);

assign xor_ln895_445_fu_35008_p2 = (p_Result_727_reg_43440 ^ 1'd1);

assign xor_ln895_446_fu_35066_p2 = (p_Result_729_reg_43460 ^ 1'd1);

assign xor_ln895_447_fu_35124_p2 = (p_Result_731_reg_43480 ^ 1'd1);

assign xor_ln895_448_fu_35182_p2 = (p_Result_733_reg_43500 ^ 1'd1);

assign xor_ln895_449_fu_35276_p2 = (p_Result_735_fu_35254_p3 ^ 1'd1);

assign xor_ln895_450_fu_35378_p2 = (p_Result_737_fu_35356_p3 ^ 1'd1);

assign xor_ln895_451_fu_35480_p2 = (p_Result_739_fu_35458_p3 ^ 1'd1);

assign xor_ln895_452_fu_35582_p2 = (p_Result_741_fu_35560_p3 ^ 1'd1);

assign xor_ln895_453_fu_35684_p2 = (p_Result_743_fu_35662_p3 ^ 1'd1);

assign xor_ln895_454_fu_35786_p2 = (p_Result_745_fu_35764_p3 ^ 1'd1);

assign xor_ln895_455_fu_35888_p2 = (p_Result_747_fu_35866_p3 ^ 1'd1);

assign xor_ln895_456_fu_35990_p2 = (p_Result_749_fu_35968_p3 ^ 1'd1);

assign xor_ln895_457_fu_36092_p2 = (p_Result_751_fu_36070_p3 ^ 1'd1);

assign xor_ln895_458_fu_36194_p2 = (p_Result_753_fu_36172_p3 ^ 1'd1);

assign xor_ln895_459_fu_36296_p2 = (p_Result_755_fu_36274_p3 ^ 1'd1);

assign xor_ln895_460_fu_36398_p2 = (p_Result_757_fu_36376_p3 ^ 1'd1);

assign xor_ln895_461_fu_36500_p2 = (p_Result_759_fu_36478_p3 ^ 1'd1);

assign xor_ln895_462_fu_36602_p2 = (p_Result_761_fu_36580_p3 ^ 1'd1);

assign xor_ln895_463_fu_36704_p2 = (p_Result_763_fu_36682_p3 ^ 1'd1);

assign xor_ln895_464_fu_36806_p2 = (p_Result_765_fu_36784_p3 ^ 1'd1);

assign xor_ln895_465_fu_36908_p2 = (p_Result_767_fu_36886_p3 ^ 1'd1);

assign xor_ln895_466_fu_37010_p2 = (p_Result_769_fu_36988_p3 ^ 1'd1);

assign xor_ln895_467_fu_39436_p2 = (p_Result_771_fu_39415_p3 ^ 1'd1);

assign xor_ln895_468_fu_39536_p2 = (p_Result_773_fu_39515_p3 ^ 1'd1);

assign xor_ln895_469_fu_39636_p2 = (p_Result_775_fu_39615_p3 ^ 1'd1);

assign xor_ln895_470_fu_39736_p2 = (p_Result_777_fu_39715_p3 ^ 1'd1);

assign xor_ln895_471_fu_39836_p2 = (p_Result_779_fu_39815_p3 ^ 1'd1);

assign xor_ln895_472_fu_39936_p2 = (p_Result_781_fu_39915_p3 ^ 1'd1);

assign xor_ln895_473_fu_40036_p2 = (p_Result_783_fu_40015_p3 ^ 1'd1);

assign xor_ln895_474_fu_40136_p2 = (p_Result_785_fu_40115_p3 ^ 1'd1);

assign xor_ln895_475_fu_40236_p2 = (p_Result_787_fu_40215_p3 ^ 1'd1);

assign xor_ln895_476_fu_40338_p2 = (p_Result_789_fu_40316_p3 ^ 1'd1);

assign xor_ln895_477_fu_40440_p2 = (p_Result_791_fu_40418_p3 ^ 1'd1);

assign xor_ln895_478_fu_40542_p2 = (p_Result_793_fu_40520_p3 ^ 1'd1);

assign xor_ln895_479_fu_40644_p2 = (p_Result_795_fu_40622_p3 ^ 1'd1);

assign xor_ln895_480_fu_40746_p2 = (p_Result_797_fu_40724_p3 ^ 1'd1);

assign xor_ln895_481_fu_40848_p2 = (p_Result_799_fu_40826_p3 ^ 1'd1);

assign xor_ln895_482_fu_40950_p2 = (p_Result_801_fu_40928_p3 ^ 1'd1);

assign xor_ln895_483_fu_41052_p2 = (p_Result_803_fu_41030_p3 ^ 1'd1);

assign xor_ln895_484_fu_41154_p2 = (p_Result_805_fu_41132_p3 ^ 1'd1);

assign xor_ln895_fu_19024_p2 = (deleted_zeros_fu_18989_p2 ^ 1'd1);

assign xor_ln896_243_fu_19046_p2 = (deleted_ones_fu_19014_p2 ^ 1'd1);

assign xor_ln896_244_fu_19094_p2 = (p_Result_407_reg_41381 ^ 1'd1);

assign xor_ln896_245_fu_19171_p2 = (deleted_ones_162_fu_19139_p2 ^ 1'd1);

assign xor_ln896_246_fu_19219_p2 = (p_Result_410_reg_41412 ^ 1'd1);

assign xor_ln896_247_fu_19296_p2 = (deleted_ones_163_fu_19264_p2 ^ 1'd1);

assign xor_ln896_248_fu_19344_p2 = (p_Result_413_reg_41443 ^ 1'd1);

assign xor_ln896_249_fu_19421_p2 = (deleted_ones_164_fu_19389_p2 ^ 1'd1);

assign xor_ln896_250_fu_19469_p2 = (p_Result_416_reg_41474 ^ 1'd1);

assign xor_ln896_251_fu_19546_p2 = (deleted_ones_165_fu_19514_p2 ^ 1'd1);

assign xor_ln896_252_fu_19594_p2 = (p_Result_419_reg_41505 ^ 1'd1);

assign xor_ln896_253_fu_19671_p2 = (deleted_ones_166_fu_19639_p2 ^ 1'd1);

assign xor_ln896_254_fu_19719_p2 = (p_Result_422_reg_41536 ^ 1'd1);

assign xor_ln896_255_fu_19796_p2 = (deleted_ones_167_fu_19764_p2 ^ 1'd1);

assign xor_ln896_256_fu_19844_p2 = (p_Result_425_reg_41567 ^ 1'd1);

assign xor_ln896_257_fu_19921_p2 = (deleted_ones_168_fu_19889_p2 ^ 1'd1);

assign xor_ln896_258_fu_19969_p2 = (p_Result_428_reg_41598 ^ 1'd1);

assign xor_ln896_259_fu_20046_p2 = (deleted_ones_169_fu_20014_p2 ^ 1'd1);

assign xor_ln896_260_fu_20115_p2 = (p_Result_431_fu_20107_p3 ^ 1'd1);

assign xor_ln896_261_fu_20195_p2 = (deleted_ones_170_fu_20162_p2 ^ 1'd1);

assign xor_ln896_262_fu_20264_p2 = (p_Result_434_fu_20256_p3 ^ 1'd1);

assign xor_ln896_263_fu_20344_p2 = (deleted_ones_171_fu_20311_p2 ^ 1'd1);

assign xor_ln896_264_fu_20413_p2 = (p_Result_437_fu_20405_p3 ^ 1'd1);

assign xor_ln896_265_fu_20493_p2 = (deleted_ones_172_fu_20460_p2 ^ 1'd1);

assign xor_ln896_266_fu_20562_p2 = (p_Result_440_fu_20554_p3 ^ 1'd1);

assign xor_ln896_267_fu_20642_p2 = (deleted_ones_173_fu_20609_p2 ^ 1'd1);

assign xor_ln896_268_fu_20711_p2 = (p_Result_443_fu_20703_p3 ^ 1'd1);

assign xor_ln896_269_fu_20791_p2 = (deleted_ones_174_fu_20758_p2 ^ 1'd1);

assign xor_ln896_270_fu_18183_p2 = (p_Result_446_fu_18175_p3 ^ 1'd1);

assign xor_ln896_271_fu_18277_p2 = (deleted_ones_175_fu_18241_p2 ^ 1'd1);

assign xor_ln896_272_fu_20877_p2 = (p_Result_449_fu_20869_p3 ^ 1'd1);

assign xor_ln896_273_fu_20957_p2 = (deleted_ones_176_fu_20924_p2 ^ 1'd1);

assign xor_ln896_274_fu_21026_p2 = (p_Result_452_fu_21018_p3 ^ 1'd1);

assign xor_ln896_275_fu_21106_p2 = (deleted_ones_177_fu_21073_p2 ^ 1'd1);

assign xor_ln896_276_fu_21175_p2 = (p_Result_455_fu_21167_p3 ^ 1'd1);

assign xor_ln896_277_fu_21255_p2 = (deleted_ones_178_fu_21222_p2 ^ 1'd1);

assign xor_ln896_278_fu_21320_p2 = (p_Result_458_fu_21312_p3 ^ 1'd1);

assign xor_ln896_279_fu_21400_p2 = (deleted_ones_179_fu_21367_p2 ^ 1'd1);

assign xor_ln896_280_fu_21465_p2 = (p_Result_461_fu_21457_p3 ^ 1'd1);

assign xor_ln896_281_fu_21545_p2 = (deleted_ones_180_fu_21512_p2 ^ 1'd1);

assign xor_ln896_282_fu_21594_p2 = (p_Result_464_fu_21586_p3 ^ 1'd1);

assign xor_ln896_283_fu_21674_p2 = (deleted_ones_181_fu_21641_p2 ^ 1'd1);

assign xor_ln896_284_fu_21719_p2 = (p_Result_467_fu_21711_p3 ^ 1'd1);

assign xor_ln896_285_fu_21799_p2 = (deleted_ones_182_fu_21766_p2 ^ 1'd1);

assign xor_ln896_286_fu_21864_p2 = (p_Result_470_fu_21856_p3 ^ 1'd1);

assign xor_ln896_287_fu_21944_p2 = (deleted_ones_183_fu_21911_p2 ^ 1'd1);

assign xor_ln896_288_fu_21993_p2 = (p_Result_473_fu_21985_p3 ^ 1'd1);

assign xor_ln896_289_fu_22073_p2 = (deleted_ones_184_fu_22040_p2 ^ 1'd1);

assign xor_ln896_290_fu_22122_p2 = (p_Result_476_fu_22114_p3 ^ 1'd1);

assign xor_ln896_291_fu_22202_p2 = (deleted_ones_185_fu_22169_p2 ^ 1'd1);

assign xor_ln896_292_fu_22251_p2 = (p_Result_479_fu_22243_p3 ^ 1'd1);

assign xor_ln896_293_fu_22331_p2 = (deleted_ones_186_fu_22298_p2 ^ 1'd1);

assign xor_ln896_294_fu_22380_p2 = (p_Result_482_fu_22372_p3 ^ 1'd1);

assign xor_ln896_295_fu_22460_p2 = (deleted_ones_187_fu_22427_p2 ^ 1'd1);

assign xor_ln896_296_fu_25544_p2 = (p_Result_485_reg_42269 ^ 1'd1);

assign xor_ln896_297_fu_25621_p2 = (deleted_ones_188_fu_25589_p2 ^ 1'd1);

assign xor_ln896_298_fu_25669_p2 = (p_Result_488_reg_42300 ^ 1'd1);

assign xor_ln896_299_fu_25746_p2 = (deleted_ones_189_fu_25714_p2 ^ 1'd1);

assign xor_ln896_300_fu_25794_p2 = (p_Result_491_reg_42331 ^ 1'd1);

assign xor_ln896_301_fu_25871_p2 = (deleted_ones_190_fu_25839_p2 ^ 1'd1);

assign xor_ln896_302_fu_25919_p2 = (p_Result_494_reg_42362 ^ 1'd1);

assign xor_ln896_303_fu_25996_p2 = (deleted_ones_191_fu_25964_p2 ^ 1'd1);

assign xor_ln896_304_fu_26044_p2 = (p_Result_497_reg_42393 ^ 1'd1);

assign xor_ln896_305_fu_26121_p2 = (deleted_ones_192_fu_26089_p2 ^ 1'd1);

assign xor_ln896_306_fu_26169_p2 = (p_Result_500_reg_42424 ^ 1'd1);

assign xor_ln896_307_fu_26246_p2 = (deleted_ones_193_fu_26214_p2 ^ 1'd1);

assign xor_ln896_308_fu_22965_p2 = (p_Result_503_fu_22957_p3 ^ 1'd1);

assign xor_ln896_309_fu_23059_p2 = (deleted_ones_194_fu_23023_p2 ^ 1'd1);

assign xor_ln896_310_fu_26311_p2 = (p_Result_506_reg_42470 ^ 1'd1);

assign xor_ln896_311_fu_26388_p2 = (deleted_ones_195_fu_26356_p2 ^ 1'd1);

assign xor_ln896_312_fu_26436_p2 = (p_Result_509_reg_42501 ^ 1'd1);

assign xor_ln896_313_fu_26513_p2 = (deleted_ones_196_fu_26481_p2 ^ 1'd1);

assign xor_ln896_314_fu_26578_p2 = (p_Result_512_fu_26570_p3 ^ 1'd1);

assign xor_ln896_315_fu_26658_p2 = (deleted_ones_197_fu_26625_p2 ^ 1'd1);

assign xor_ln896_316_fu_26727_p2 = (p_Result_515_fu_26719_p3 ^ 1'd1);

assign xor_ln896_317_fu_26807_p2 = (deleted_ones_198_fu_26774_p2 ^ 1'd1);

assign xor_ln896_318_fu_26876_p2 = (p_Result_518_fu_26868_p3 ^ 1'd1);

assign xor_ln896_319_fu_26956_p2 = (deleted_ones_199_fu_26923_p2 ^ 1'd1);

assign xor_ln896_320_fu_27025_p2 = (p_Result_521_fu_27017_p3 ^ 1'd1);

assign xor_ln896_321_fu_27105_p2 = (deleted_ones_200_fu_27072_p2 ^ 1'd1);

assign xor_ln896_322_fu_27174_p2 = (p_Result_524_fu_27166_p3 ^ 1'd1);

assign xor_ln896_323_fu_27254_p2 = (deleted_ones_201_fu_27221_p2 ^ 1'd1);

assign xor_ln896_324_fu_27323_p2 = (p_Result_527_fu_27315_p3 ^ 1'd1);

assign xor_ln896_325_fu_27403_p2 = (deleted_ones_202_fu_27370_p2 ^ 1'd1);

assign xor_ln896_326_fu_27472_p2 = (p_Result_530_fu_27464_p3 ^ 1'd1);

assign xor_ln896_327_fu_27552_p2 = (deleted_ones_203_fu_27519_p2 ^ 1'd1);

assign xor_ln896_328_fu_27621_p2 = (p_Result_533_fu_27613_p3 ^ 1'd1);

assign xor_ln896_329_fu_27701_p2 = (deleted_ones_204_fu_27668_p2 ^ 1'd1);

assign xor_ln896_330_fu_27770_p2 = (p_Result_536_fu_27762_p3 ^ 1'd1);

assign xor_ln896_331_fu_27850_p2 = (deleted_ones_205_fu_27817_p2 ^ 1'd1);

assign xor_ln896_332_fu_27993_p2 = (p_Result_539_fu_27985_p3 ^ 1'd1);

assign xor_ln896_333_fu_28087_p2 = (deleted_ones_206_fu_28051_p2 ^ 1'd1);

assign xor_ln896_334_fu_31342_p2 = (p_Result_542_reg_42862 ^ 1'd1);

assign xor_ln896_335_fu_31419_p2 = (deleted_ones_207_fu_31387_p2 ^ 1'd1);

assign xor_ln896_336_fu_31467_p2 = (p_Result_545_reg_42893 ^ 1'd1);

assign xor_ln896_337_fu_31544_p2 = (deleted_ones_208_fu_31512_p2 ^ 1'd1);

assign xor_ln896_338_fu_31592_p2 = (p_Result_548_reg_42924 ^ 1'd1);

assign xor_ln896_339_fu_31669_p2 = (deleted_ones_209_fu_31637_p2 ^ 1'd1);

assign xor_ln896_340_fu_31717_p2 = (p_Result_551_reg_42955 ^ 1'd1);

assign xor_ln896_341_fu_31794_p2 = (deleted_ones_210_fu_31762_p2 ^ 1'd1);

assign xor_ln896_342_fu_31842_p2 = (p_Result_554_reg_42986 ^ 1'd1);

assign xor_ln896_343_fu_31919_p2 = (deleted_ones_211_fu_31887_p2 ^ 1'd1);

assign xor_ln896_344_fu_31967_p2 = (p_Result_557_reg_43017 ^ 1'd1);

assign xor_ln896_345_fu_32044_p2 = (deleted_ones_212_fu_32012_p2 ^ 1'd1);

assign xor_ln896_346_fu_32092_p2 = (p_Result_560_reg_43048 ^ 1'd1);

assign xor_ln896_347_fu_32169_p2 = (deleted_ones_213_fu_32137_p2 ^ 1'd1);

assign xor_ln896_348_fu_32217_p2 = (p_Result_563_reg_43079 ^ 1'd1);

assign xor_ln896_349_fu_32294_p2 = (deleted_ones_214_fu_32262_p2 ^ 1'd1);

assign xor_ln896_350_fu_32363_p2 = (p_Result_566_fu_32355_p3 ^ 1'd1);

assign xor_ln896_351_fu_32443_p2 = (deleted_ones_215_fu_32410_p2 ^ 1'd1);

assign xor_ln896_352_fu_32512_p2 = (p_Result_569_fu_32504_p3 ^ 1'd1);

assign xor_ln896_353_fu_32592_p2 = (deleted_ones_216_fu_32559_p2 ^ 1'd1);

assign xor_ln896_354_fu_32661_p2 = (p_Result_572_fu_32653_p3 ^ 1'd1);

assign xor_ln896_355_fu_32741_p2 = (deleted_ones_217_fu_32708_p2 ^ 1'd1);

assign xor_ln896_356_fu_32810_p2 = (p_Result_575_fu_32802_p3 ^ 1'd1);

assign xor_ln896_357_fu_32890_p2 = (deleted_ones_218_fu_32857_p2 ^ 1'd1);

assign xor_ln896_358_fu_32959_p2 = (p_Result_578_fu_32951_p3 ^ 1'd1);

assign xor_ln896_359_fu_33039_p2 = (deleted_ones_219_fu_33006_p2 ^ 1'd1);

assign xor_ln896_360_fu_33108_p2 = (p_Result_581_fu_33100_p3 ^ 1'd1);

assign xor_ln896_361_fu_33188_p2 = (deleted_ones_220_fu_33155_p2 ^ 1'd1);

assign xor_ln896_362_fu_33257_p2 = (p_Result_584_fu_33249_p3 ^ 1'd1);

assign xor_ln896_363_fu_33337_p2 = (deleted_ones_221_fu_33304_p2 ^ 1'd1);

assign xor_ln896_364_fu_33406_p2 = (p_Result_587_fu_33398_p3 ^ 1'd1);

assign xor_ln896_365_fu_33486_p2 = (deleted_ones_222_fu_33453_p2 ^ 1'd1);

assign xor_ln896_366_fu_29060_p2 = (p_Result_590_fu_29052_p3 ^ 1'd1);

assign xor_ln896_367_fu_29154_p2 = (deleted_ones_223_fu_29118_p2 ^ 1'd1);

assign xor_ln896_368_fu_37076_p2 = (p_Result_593_reg_43537 ^ 1'd1);

assign xor_ln896_369_fu_37153_p2 = (deleted_ones_224_fu_37121_p2 ^ 1'd1);

assign xor_ln896_370_fu_37200_p2 = (p_Result_596_reg_43568 ^ 1'd1);

assign xor_ln896_371_fu_37277_p2 = (deleted_ones_225_fu_37245_p2 ^ 1'd1);

assign xor_ln896_372_fu_37325_p2 = (p_Result_599_reg_43599 ^ 1'd1);

assign xor_ln896_373_fu_37402_p2 = (deleted_ones_226_fu_37370_p2 ^ 1'd1);

assign xor_ln896_374_fu_37450_p2 = (p_Result_602_reg_43630 ^ 1'd1);

assign xor_ln896_375_fu_37527_p2 = (deleted_ones_227_fu_37495_p2 ^ 1'd1);

assign xor_ln896_376_fu_37575_p2 = (p_Result_605_reg_43661 ^ 1'd1);

assign xor_ln896_377_fu_37652_p2 = (deleted_ones_228_fu_37620_p2 ^ 1'd1);

assign xor_ln896_378_fu_37700_p2 = (p_Result_608_reg_43692 ^ 1'd1);

assign xor_ln896_379_fu_37777_p2 = (deleted_ones_229_fu_37745_p2 ^ 1'd1);

assign xor_ln896_380_fu_37825_p2 = (p_Result_611_reg_43723 ^ 1'd1);

assign xor_ln896_381_fu_37902_p2 = (deleted_ones_230_fu_37870_p2 ^ 1'd1);

assign xor_ln896_382_fu_37950_p2 = (p_Result_614_reg_43754 ^ 1'd1);

assign xor_ln896_383_fu_38027_p2 = (deleted_ones_231_fu_37995_p2 ^ 1'd1);

assign xor_ln896_384_fu_38075_p2 = (p_Result_617_reg_43785 ^ 1'd1);

assign xor_ln896_385_fu_38152_p2 = (deleted_ones_232_fu_38120_p2 ^ 1'd1);

assign xor_ln896_386_fu_38217_p2 = (p_Result_620_fu_38209_p3 ^ 1'd1);

assign xor_ln896_387_fu_38297_p2 = (deleted_ones_233_fu_38264_p2 ^ 1'd1);

assign xor_ln896_388_fu_38366_p2 = (p_Result_623_fu_38358_p3 ^ 1'd1);

assign xor_ln896_389_fu_38446_p2 = (deleted_ones_234_fu_38413_p2 ^ 1'd1);

assign xor_ln896_390_fu_38515_p2 = (p_Result_626_fu_38507_p3 ^ 1'd1);

assign xor_ln896_391_fu_38595_p2 = (deleted_ones_235_fu_38562_p2 ^ 1'd1);

assign xor_ln896_392_fu_38664_p2 = (p_Result_629_fu_38656_p3 ^ 1'd1);

assign xor_ln896_393_fu_38744_p2 = (deleted_ones_236_fu_38711_p2 ^ 1'd1);

assign xor_ln896_394_fu_38813_p2 = (p_Result_632_fu_38805_p3 ^ 1'd1);

assign xor_ln896_395_fu_38893_p2 = (deleted_ones_237_fu_38860_p2 ^ 1'd1);

assign xor_ln896_396_fu_38962_p2 = (p_Result_635_fu_38954_p3 ^ 1'd1);

assign xor_ln896_397_fu_39042_p2 = (deleted_ones_238_fu_39009_p2 ^ 1'd1);

assign xor_ln896_398_fu_39111_p2 = (p_Result_638_fu_39103_p3 ^ 1'd1);

assign xor_ln896_399_fu_39191_p2 = (deleted_ones_239_fu_39158_p2 ^ 1'd1);

assign xor_ln896_400_fu_34552_p2 = (p_Result_641_fu_34544_p3 ^ 1'd1);

assign xor_ln896_401_fu_34646_p2 = (deleted_ones_240_fu_34610_p2 ^ 1'd1);

assign xor_ln896_402_fu_39277_p2 = (p_Result_644_fu_39269_p3 ^ 1'd1);

assign xor_ln896_403_fu_39357_p2 = (deleted_ones_241_fu_39324_p2 ^ 1'd1);

assign xor_ln896_404_fu_23666_p2 = (p_Result_646_fu_23646_p3 ^ 1'd1);

assign xor_ln896_405_fu_23764_p2 = (p_Result_648_fu_23744_p3 ^ 1'd1);

assign xor_ln896_406_fu_23862_p2 = (p_Result_650_fu_23842_p3 ^ 1'd1);

assign xor_ln896_407_fu_23960_p2 = (p_Result_652_fu_23940_p3 ^ 1'd1);

assign xor_ln896_408_fu_24058_p2 = (p_Result_654_fu_24038_p3 ^ 1'd1);

assign xor_ln896_409_fu_24156_p2 = (p_Result_656_fu_24136_p3 ^ 1'd1);

assign xor_ln896_410_fu_24254_p2 = (p_Result_658_fu_24234_p3 ^ 1'd1);

assign xor_ln896_411_fu_24352_p2 = (p_Result_660_fu_24332_p3 ^ 1'd1);

assign xor_ln896_412_fu_24450_p2 = (p_Result_662_fu_24430_p3 ^ 1'd1);

assign xor_ln896_413_fu_24552_p2 = (p_Result_664_fu_24532_p3 ^ 1'd1);

assign xor_ln896_414_fu_24654_p2 = (p_Result_666_fu_24634_p3 ^ 1'd1);

assign xor_ln896_415_fu_24756_p2 = (p_Result_668_fu_24736_p3 ^ 1'd1);

assign xor_ln896_416_fu_24858_p2 = (p_Result_670_fu_24838_p3 ^ 1'd1);

assign xor_ln896_417_fu_24960_p2 = (p_Result_672_fu_24940_p3 ^ 1'd1);

assign xor_ln896_418_fu_25062_p2 = (p_Result_674_fu_25042_p3 ^ 1'd1);

assign xor_ln896_419_fu_25164_p2 = (p_Result_676_fu_25144_p3 ^ 1'd1);

assign xor_ln896_420_fu_25266_p2 = (p_Result_678_fu_25246_p3 ^ 1'd1);

assign xor_ln896_421_fu_25368_p2 = (p_Result_680_fu_25348_p3 ^ 1'd1);

assign xor_ln896_422_fu_29228_p2 = (p_Result_682_fu_29208_p3 ^ 1'd1);

assign xor_ln896_423_fu_29328_p2 = (p_Result_684_fu_29308_p3 ^ 1'd1);

assign xor_ln896_424_fu_29428_p2 = (p_Result_686_fu_29408_p3 ^ 1'd1);

assign xor_ln896_425_fu_29526_p2 = (p_Result_688_fu_29506_p3 ^ 1'd1);

assign xor_ln896_426_fu_29626_p2 = (p_Result_690_fu_29606_p3 ^ 1'd1);

assign xor_ln896_427_fu_29726_p2 = (p_Result_692_fu_29706_p3 ^ 1'd1);

assign xor_ln896_428_fu_29826_p2 = (p_Result_694_fu_29806_p3 ^ 1'd1);

assign xor_ln896_429_fu_29926_p2 = (p_Result_696_fu_29906_p3 ^ 1'd1);

assign xor_ln896_430_fu_30026_p2 = (p_Result_698_fu_30006_p3 ^ 1'd1);

assign xor_ln896_431_fu_30128_p2 = (p_Result_700_fu_30108_p3 ^ 1'd1);

assign xor_ln896_432_fu_30230_p2 = (p_Result_702_fu_30210_p3 ^ 1'd1);

assign xor_ln896_433_fu_30332_p2 = (p_Result_704_fu_30312_p3 ^ 1'd1);

assign xor_ln896_434_fu_30434_p2 = (p_Result_706_fu_30414_p3 ^ 1'd1);

assign xor_ln896_435_fu_30536_p2 = (p_Result_708_fu_30516_p3 ^ 1'd1);

assign xor_ln896_436_fu_30638_p2 = (p_Result_710_fu_30618_p3 ^ 1'd1);

assign xor_ln896_437_fu_30740_p2 = (p_Result_712_fu_30720_p3 ^ 1'd1);

assign xor_ln896_438_fu_30842_p2 = (p_Result_714_fu_30822_p3 ^ 1'd1);

assign xor_ln896_439_fu_30944_p2 = (p_Result_716_fu_30924_p3 ^ 1'd1);

assign xor_ln896_440_fu_34728_p2 = (p_Result_718_reg_43353 ^ 1'd1);

assign xor_ln896_441_fu_34786_p2 = (p_Result_720_reg_43373 ^ 1'd1);

assign xor_ln896_442_fu_34844_p2 = (p_Result_722_reg_43393 ^ 1'd1);

assign xor_ln896_443_fu_34902_p2 = (p_Result_724_reg_43413 ^ 1'd1);

assign xor_ln896_444_fu_34960_p2 = (p_Result_726_reg_43433 ^ 1'd1);

assign xor_ln896_445_fu_35018_p2 = (p_Result_728_reg_43453 ^ 1'd1);

assign xor_ln896_446_fu_35076_p2 = (p_Result_730_reg_43473 ^ 1'd1);

assign xor_ln896_447_fu_35134_p2 = (p_Result_732_reg_43493 ^ 1'd1);

assign xor_ln896_448_fu_35192_p2 = (p_Result_734_reg_43513 ^ 1'd1);

assign xor_ln896_449_fu_35288_p2 = (p_Result_736_fu_35268_p3 ^ 1'd1);

assign xor_ln896_450_fu_35390_p2 = (p_Result_738_fu_35370_p3 ^ 1'd1);

assign xor_ln896_451_fu_35492_p2 = (p_Result_740_fu_35472_p3 ^ 1'd1);

assign xor_ln896_452_fu_35594_p2 = (p_Result_742_fu_35574_p3 ^ 1'd1);

assign xor_ln896_453_fu_35696_p2 = (p_Result_744_fu_35676_p3 ^ 1'd1);

assign xor_ln896_454_fu_35798_p2 = (p_Result_746_fu_35778_p3 ^ 1'd1);

assign xor_ln896_455_fu_35900_p2 = (p_Result_748_fu_35880_p3 ^ 1'd1);

assign xor_ln896_456_fu_36002_p2 = (p_Result_750_fu_35982_p3 ^ 1'd1);

assign xor_ln896_457_fu_36104_p2 = (p_Result_752_fu_36084_p3 ^ 1'd1);

assign xor_ln896_458_fu_36206_p2 = (p_Result_754_fu_36186_p3 ^ 1'd1);

assign xor_ln896_459_fu_36308_p2 = (p_Result_756_fu_36288_p3 ^ 1'd1);

assign xor_ln896_460_fu_36410_p2 = (p_Result_758_fu_36390_p3 ^ 1'd1);

assign xor_ln896_461_fu_36512_p2 = (p_Result_760_fu_36492_p3 ^ 1'd1);

assign xor_ln896_462_fu_36614_p2 = (p_Result_762_fu_36594_p3 ^ 1'd1);

assign xor_ln896_463_fu_36716_p2 = (p_Result_764_fu_36696_p3 ^ 1'd1);

assign xor_ln896_464_fu_36818_p2 = (p_Result_766_fu_36798_p3 ^ 1'd1);

assign xor_ln896_465_fu_36920_p2 = (p_Result_768_fu_36900_p3 ^ 1'd1);

assign xor_ln896_466_fu_37022_p2 = (p_Result_770_fu_37002_p3 ^ 1'd1);

assign xor_ln896_467_fu_39448_p2 = (p_Result_772_fu_39428_p3 ^ 1'd1);

assign xor_ln896_468_fu_39548_p2 = (p_Result_774_fu_39528_p3 ^ 1'd1);

assign xor_ln896_469_fu_39648_p2 = (p_Result_776_fu_39628_p3 ^ 1'd1);

assign xor_ln896_470_fu_39748_p2 = (p_Result_778_fu_39728_p3 ^ 1'd1);

assign xor_ln896_471_fu_39848_p2 = (p_Result_780_fu_39828_p3 ^ 1'd1);

assign xor_ln896_472_fu_39948_p2 = (p_Result_782_fu_39928_p3 ^ 1'd1);

assign xor_ln896_473_fu_40048_p2 = (p_Result_784_fu_40028_p3 ^ 1'd1);

assign xor_ln896_474_fu_40148_p2 = (p_Result_786_fu_40128_p3 ^ 1'd1);

assign xor_ln896_475_fu_40248_p2 = (p_Result_788_fu_40228_p3 ^ 1'd1);

assign xor_ln896_476_fu_40350_p2 = (p_Result_790_fu_40330_p3 ^ 1'd1);

assign xor_ln896_477_fu_40452_p2 = (p_Result_792_fu_40432_p3 ^ 1'd1);

assign xor_ln896_478_fu_40554_p2 = (p_Result_794_fu_40534_p3 ^ 1'd1);

assign xor_ln896_479_fu_40656_p2 = (p_Result_796_fu_40636_p3 ^ 1'd1);

assign xor_ln896_480_fu_40758_p2 = (p_Result_798_fu_40738_p3 ^ 1'd1);

assign xor_ln896_481_fu_40860_p2 = (p_Result_800_fu_40840_p3 ^ 1'd1);

assign xor_ln896_482_fu_40962_p2 = (p_Result_802_fu_40942_p3 ^ 1'd1);

assign xor_ln896_483_fu_41064_p2 = (p_Result_804_fu_41044_p3 ^ 1'd1);

assign xor_ln896_484_fu_41166_p2 = (p_Result_806_fu_41146_p3 ^ 1'd1);

assign xor_ln896_485_fu_19058_p2 = (or_ln896_fu_19052_p2 ^ and_ln891_fu_19019_p2);

assign xor_ln896_486_fu_19183_p2 = (or_ln896_81_fu_19177_p2 ^ and_ln891_81_fu_19144_p2);

assign xor_ln896_487_fu_19308_p2 = (or_ln896_82_fu_19302_p2 ^ and_ln891_82_fu_19269_p2);

assign xor_ln896_488_fu_19433_p2 = (or_ln896_83_fu_19427_p2 ^ and_ln891_83_fu_19394_p2);

assign xor_ln896_489_fu_19558_p2 = (or_ln896_84_fu_19552_p2 ^ and_ln891_84_fu_19519_p2);

assign xor_ln896_490_fu_19683_p2 = (or_ln896_85_fu_19677_p2 ^ and_ln891_85_fu_19644_p2);

assign xor_ln896_491_fu_19808_p2 = (or_ln896_86_fu_19802_p2 ^ and_ln891_86_fu_19769_p2);

assign xor_ln896_492_fu_19933_p2 = (or_ln896_87_fu_19927_p2 ^ and_ln891_87_fu_19894_p2);

assign xor_ln896_493_fu_20058_p2 = (or_ln896_88_fu_20052_p2 ^ and_ln891_88_fu_20019_p2);

assign xor_ln896_494_fu_20207_p2 = (or_ln896_89_fu_20201_p2 ^ and_ln891_89_fu_20167_p2);

assign xor_ln896_495_fu_20356_p2 = (or_ln896_90_fu_20350_p2 ^ and_ln891_90_fu_20316_p2);

assign xor_ln896_496_fu_20505_p2 = (or_ln896_91_fu_20499_p2 ^ and_ln891_91_fu_20465_p2);

assign xor_ln896_497_fu_20654_p2 = (or_ln896_92_fu_20648_p2 ^ and_ln891_92_fu_20614_p2);

assign xor_ln896_498_fu_20803_p2 = (or_ln896_93_fu_20797_p2 ^ and_ln891_93_fu_20763_p2);

assign xor_ln896_499_fu_18289_p2 = (or_ln896_94_fu_18283_p2 ^ and_ln891_94_fu_18247_p2);

assign xor_ln896_500_fu_20969_p2 = (or_ln896_95_fu_20963_p2 ^ and_ln891_95_fu_20929_p2);

assign xor_ln896_501_fu_21118_p2 = (or_ln896_96_fu_21112_p2 ^ and_ln891_96_fu_21078_p2);

assign xor_ln896_502_fu_21267_p2 = (or_ln896_97_fu_21261_p2 ^ and_ln891_97_fu_21227_p2);

assign xor_ln896_503_fu_21412_p2 = (or_ln896_98_fu_21406_p2 ^ and_ln891_98_fu_21372_p2);

assign xor_ln896_504_fu_21557_p2 = (or_ln896_99_fu_21551_p2 ^ and_ln891_99_fu_21517_p2);

assign xor_ln896_505_fu_21686_p2 = (or_ln896_100_fu_21680_p2 ^ and_ln891_100_fu_21646_p2);

assign xor_ln896_506_fu_21811_p2 = (or_ln896_101_fu_21805_p2 ^ and_ln891_101_fu_21771_p2);

assign xor_ln896_507_fu_21956_p2 = (or_ln896_102_fu_21950_p2 ^ and_ln891_102_fu_21916_p2);

assign xor_ln896_508_fu_22085_p2 = (or_ln896_103_fu_22079_p2 ^ and_ln891_103_fu_22045_p2);

assign xor_ln896_509_fu_22214_p2 = (or_ln896_104_fu_22208_p2 ^ and_ln891_104_fu_22174_p2);

assign xor_ln896_510_fu_22343_p2 = (or_ln896_105_fu_22337_p2 ^ and_ln891_105_fu_22303_p2);

assign xor_ln896_511_fu_22472_p2 = (or_ln896_106_fu_22466_p2 ^ and_ln891_106_fu_22432_p2);

assign xor_ln896_512_fu_25633_p2 = (or_ln896_107_fu_25627_p2 ^ and_ln891_107_fu_25594_p2);

assign xor_ln896_513_fu_25758_p2 = (or_ln896_108_fu_25752_p2 ^ and_ln891_108_fu_25719_p2);

assign xor_ln896_514_fu_25883_p2 = (or_ln896_109_fu_25877_p2 ^ and_ln891_109_fu_25844_p2);

assign xor_ln896_515_fu_26008_p2 = (or_ln896_110_fu_26002_p2 ^ and_ln891_110_fu_25969_p2);

assign xor_ln896_516_fu_26133_p2 = (or_ln896_111_fu_26127_p2 ^ and_ln891_111_fu_26094_p2);

assign xor_ln896_517_fu_26258_p2 = (or_ln896_112_fu_26252_p2 ^ and_ln891_112_fu_26219_p2);

assign xor_ln896_518_fu_23071_p2 = (or_ln896_113_fu_23065_p2 ^ and_ln891_113_fu_23029_p2);

assign xor_ln896_519_fu_26400_p2 = (or_ln896_114_fu_26394_p2 ^ and_ln891_114_fu_26361_p2);

assign xor_ln896_520_fu_26525_p2 = (or_ln896_115_fu_26519_p2 ^ and_ln891_115_fu_26486_p2);

assign xor_ln896_521_fu_26670_p2 = (or_ln896_116_fu_26664_p2 ^ and_ln891_116_fu_26630_p2);

assign xor_ln896_522_fu_26819_p2 = (or_ln896_117_fu_26813_p2 ^ and_ln891_117_fu_26779_p2);

assign xor_ln896_523_fu_26968_p2 = (or_ln896_118_fu_26962_p2 ^ and_ln891_118_fu_26928_p2);

assign xor_ln896_524_fu_27117_p2 = (or_ln896_119_fu_27111_p2 ^ and_ln891_119_fu_27077_p2);

assign xor_ln896_525_fu_27266_p2 = (or_ln896_120_fu_27260_p2 ^ and_ln891_120_fu_27226_p2);

assign xor_ln896_526_fu_27415_p2 = (or_ln896_121_fu_27409_p2 ^ and_ln891_121_fu_27375_p2);

assign xor_ln896_527_fu_27564_p2 = (or_ln896_122_fu_27558_p2 ^ and_ln891_122_fu_27524_p2);

assign xor_ln896_528_fu_27713_p2 = (or_ln896_123_fu_27707_p2 ^ and_ln891_123_fu_27673_p2);

assign xor_ln896_529_fu_27862_p2 = (or_ln896_124_fu_27856_p2 ^ and_ln891_124_fu_27822_p2);

assign xor_ln896_530_fu_28099_p2 = (or_ln896_125_fu_28093_p2 ^ and_ln891_125_fu_28057_p2);

assign xor_ln896_531_fu_31431_p2 = (or_ln896_126_fu_31425_p2 ^ and_ln891_126_fu_31392_p2);

assign xor_ln896_532_fu_31556_p2 = (or_ln896_127_fu_31550_p2 ^ and_ln891_127_fu_31517_p2);

assign xor_ln896_533_fu_31681_p2 = (or_ln896_128_fu_31675_p2 ^ and_ln891_128_fu_31642_p2);

assign xor_ln896_534_fu_31806_p2 = (or_ln896_129_fu_31800_p2 ^ and_ln891_129_fu_31767_p2);

assign xor_ln896_535_fu_31931_p2 = (or_ln896_130_fu_31925_p2 ^ and_ln891_130_fu_31892_p2);

assign xor_ln896_536_fu_32056_p2 = (or_ln896_131_fu_32050_p2 ^ and_ln891_131_fu_32017_p2);

assign xor_ln896_537_fu_32181_p2 = (or_ln896_132_fu_32175_p2 ^ and_ln891_132_fu_32142_p2);

assign xor_ln896_538_fu_32306_p2 = (or_ln896_133_fu_32300_p2 ^ and_ln891_133_fu_32267_p2);

assign xor_ln896_539_fu_32455_p2 = (or_ln896_134_fu_32449_p2 ^ and_ln891_134_fu_32415_p2);

assign xor_ln896_540_fu_32604_p2 = (or_ln896_135_fu_32598_p2 ^ and_ln891_135_fu_32564_p2);

assign xor_ln896_541_fu_32753_p2 = (or_ln896_136_fu_32747_p2 ^ and_ln891_136_fu_32713_p2);

assign xor_ln896_542_fu_32902_p2 = (or_ln896_137_fu_32896_p2 ^ and_ln891_137_fu_32862_p2);

assign xor_ln896_543_fu_33051_p2 = (or_ln896_138_fu_33045_p2 ^ and_ln891_138_fu_33011_p2);

assign xor_ln896_544_fu_33200_p2 = (or_ln896_139_fu_33194_p2 ^ and_ln891_139_fu_33160_p2);

assign xor_ln896_545_fu_33349_p2 = (or_ln896_140_fu_33343_p2 ^ and_ln891_140_fu_33309_p2);

assign xor_ln896_546_fu_33498_p2 = (or_ln896_141_fu_33492_p2 ^ and_ln891_141_fu_33458_p2);

assign xor_ln896_547_fu_29166_p2 = (or_ln896_142_fu_29160_p2 ^ and_ln891_142_fu_29124_p2);

assign xor_ln896_548_fu_37165_p2 = (or_ln896_143_fu_37159_p2 ^ and_ln891_143_fu_37126_p2);

assign xor_ln896_549_fu_37289_p2 = (or_ln896_144_fu_37283_p2 ^ and_ln891_144_fu_37250_p2);

assign xor_ln896_550_fu_37414_p2 = (or_ln896_145_fu_37408_p2 ^ and_ln891_145_fu_37375_p2);

assign xor_ln896_551_fu_37539_p2 = (or_ln896_146_fu_37533_p2 ^ and_ln891_146_fu_37500_p2);

assign xor_ln896_552_fu_37664_p2 = (or_ln896_147_fu_37658_p2 ^ and_ln891_147_fu_37625_p2);

assign xor_ln896_553_fu_37789_p2 = (or_ln896_148_fu_37783_p2 ^ and_ln891_148_fu_37750_p2);

assign xor_ln896_554_fu_37914_p2 = (or_ln896_149_fu_37908_p2 ^ and_ln891_149_fu_37875_p2);

assign xor_ln896_555_fu_38039_p2 = (or_ln896_150_fu_38033_p2 ^ and_ln891_150_fu_38000_p2);

assign xor_ln896_556_fu_38164_p2 = (or_ln896_151_fu_38158_p2 ^ and_ln891_151_fu_38125_p2);

assign xor_ln896_557_fu_38309_p2 = (or_ln896_152_fu_38303_p2 ^ and_ln891_152_fu_38269_p2);

assign xor_ln896_558_fu_38458_p2 = (or_ln896_153_fu_38452_p2 ^ and_ln891_153_fu_38418_p2);

assign xor_ln896_559_fu_38607_p2 = (or_ln896_154_fu_38601_p2 ^ and_ln891_154_fu_38567_p2);

assign xor_ln896_560_fu_38756_p2 = (or_ln896_155_fu_38750_p2 ^ and_ln891_155_fu_38716_p2);

assign xor_ln896_561_fu_38905_p2 = (or_ln896_156_fu_38899_p2 ^ and_ln891_156_fu_38865_p2);

assign xor_ln896_562_fu_39054_p2 = (or_ln896_157_fu_39048_p2 ^ and_ln891_157_fu_39014_p2);

assign xor_ln896_563_fu_39203_p2 = (or_ln896_158_fu_39197_p2 ^ and_ln891_158_fu_39163_p2);

assign xor_ln896_564_fu_34658_p2 = (or_ln896_159_fu_34652_p2 ^ and_ln891_159_fu_34616_p2);

assign xor_ln896_565_fu_39369_p2 = (or_ln896_160_fu_39363_p2 ^ and_ln891_160_fu_39329_p2);

assign xor_ln896_fu_18969_p2 = (p_Result_404_reg_41350 ^ 1'd1);

assign zext_ln377_100_fu_21577_p1 = tmp_759_reg_41934;

assign zext_ln377_101_fu_21703_p1 = tmp_765_reg_41963;

assign zext_ln377_102_fu_21847_p1 = tmp_771_reg_41992;

assign zext_ln377_103_fu_21976_p1 = tmp_777_reg_42021;

assign zext_ln377_104_fu_22105_p1 = tmp_783_reg_42050;

assign zext_ln377_105_fu_22234_p1 = tmp_789_reg_42079;

assign zext_ln377_106_fu_22363_p1 = tmp_795_reg_42108;

assign zext_ln377_107_fu_22544_p1 = tmp_801_fu_22536_p3;

assign zext_ln377_108_fu_22608_p1 = tmp_807_fu_22600_p3;

assign zext_ln377_109_fu_22672_p1 = tmp_813_fu_22664_p3;

assign zext_ln377_110_fu_22736_p1 = tmp_819_fu_22728_p3;

assign zext_ln377_111_fu_22800_p1 = tmp_825_fu_22792_p3;

assign zext_ln377_112_fu_22864_p1 = tmp_831_fu_22856_p3;

assign zext_ln377_113_fu_22948_p1 = tmp_837_reg_42120;

assign zext_ln377_114_fu_23127_p1 = tmp_843_fu_23119_p3;

assign zext_ln377_115_fu_23191_p1 = tmp_849_fu_23183_p3;

assign zext_ln377_116_fu_26561_p1 = tmp_855_reg_42532;

assign zext_ln377_117_fu_26706_p1 = tmp_861_reg_42561;

assign zext_ln377_118_fu_26855_p1 = tmp_867_reg_42590;

assign zext_ln377_119_fu_27004_p1 = tmp_873_reg_42619;

assign zext_ln377_120_fu_27153_p1 = tmp_879_reg_42648;

assign zext_ln377_121_fu_27302_p1 = tmp_885_reg_42677;

assign zext_ln377_122_fu_27451_p1 = tmp_891_reg_42706;

assign zext_ln377_123_fu_27600_p1 = tmp_897_reg_42735;

assign zext_ln377_124_fu_27749_p1 = tmp_903_reg_42764;

assign zext_ln377_125_fu_27976_p1 = tmp_909_reg_42125_pp0_iter1_reg;

assign zext_ln377_126_fu_28155_p1 = tmp_915_fu_28147_p3;

assign zext_ln377_127_fu_28219_p1 = tmp_921_fu_28211_p3;

assign zext_ln377_128_fu_28283_p1 = tmp_927_fu_28275_p3;

assign zext_ln377_129_fu_28347_p1 = tmp_933_fu_28339_p3;

assign zext_ln377_130_fu_28411_p1 = tmp_939_fu_28403_p3;

assign zext_ln377_131_fu_28475_p1 = tmp_945_fu_28467_p3;

assign zext_ln377_132_fu_28539_p1 = tmp_951_fu_28531_p3;

assign zext_ln377_133_fu_28603_p1 = tmp_957_fu_28595_p3;

assign zext_ln377_134_fu_32342_p1 = tmp_963_reg_43110;

assign zext_ln377_135_fu_32491_p1 = tmp_969_reg_43139;

assign zext_ln377_136_fu_32640_p1 = tmp_975_reg_43168;

assign zext_ln377_137_fu_32789_p1 = tmp_981_reg_43197;

assign zext_ln377_138_fu_32938_p1 = tmp_987_reg_43226;

assign zext_ln377_139_fu_33087_p1 = tmp_993_reg_43255;

assign zext_ln377_140_fu_33236_p1 = tmp_999_reg_43284;

assign zext_ln377_141_fu_33385_p1 = tmp_1005_reg_43313;

assign zext_ln377_142_fu_29043_p1 = tmp_1011_reg_42130_pp0_iter1_reg;

assign zext_ln377_143_fu_33610_p1 = tmp_1017_fu_33602_p3;

assign zext_ln377_144_fu_33674_p1 = tmp_1023_fu_33666_p3;

assign zext_ln377_145_fu_33738_p1 = tmp_1029_fu_33730_p3;

assign zext_ln377_146_fu_33802_p1 = tmp_1035_fu_33794_p3;

assign zext_ln377_147_fu_33866_p1 = tmp_1041_fu_33858_p3;

assign zext_ln377_148_fu_33930_p1 = tmp_1047_fu_33922_p3;

assign zext_ln377_149_fu_33994_p1 = tmp_1053_fu_33986_p3;

assign zext_ln377_150_fu_34058_p1 = tmp_1059_fu_34050_p3;

assign zext_ln377_151_fu_34122_p1 = tmp_1065_fu_34114_p3;

assign zext_ln377_152_fu_38200_p1 = tmp_1071_reg_43816;

assign zext_ln377_153_fu_38345_p1 = tmp_1077_reg_43845;

assign zext_ln377_154_fu_38494_p1 = tmp_1083_reg_43874;

assign zext_ln377_155_fu_38643_p1 = tmp_1089_reg_43903;

assign zext_ln377_156_fu_38792_p1 = tmp_1095_reg_43932;

assign zext_ln377_157_fu_38941_p1 = tmp_1101_reg_43961;

assign zext_ln377_158_fu_39090_p1 = tmp_1107_reg_43990;

assign zext_ln377_159_fu_34534_p1 = tmp_1113_fu_34526_p3;

assign zext_ln377_160_fu_39256_p1 = tmp_1119_reg_44034;

assign zext_ln377_81_fu_17375_p1 = tmp_645_fu_17367_p3;

assign zext_ln377_82_fu_17439_p1 = tmp_651_fu_17431_p3;

assign zext_ln377_83_fu_17503_p1 = tmp_657_fu_17495_p3;

assign zext_ln377_84_fu_17567_p1 = tmp_663_fu_17559_p3;

assign zext_ln377_85_fu_17631_p1 = tmp_669_fu_17623_p3;

assign zext_ln377_86_fu_17695_p1 = tmp_675_fu_17687_p3;

assign zext_ln377_87_fu_17759_p1 = tmp_681_fu_17751_p3;

assign zext_ln377_88_fu_17823_p1 = tmp_687_fu_17815_p3;

assign zext_ln377_89_fu_20094_p1 = tmp_693_reg_41629;

assign zext_ln377_90_fu_20243_p1 = tmp_699_reg_41658;

assign zext_ln377_91_fu_20392_p1 = tmp_705_reg_41687;

assign zext_ln377_92_fu_20541_p1 = tmp_711_reg_41716;

assign zext_ln377_93_fu_20690_p1 = tmp_717_reg_41745;

assign zext_ln377_94_fu_18165_p1 = tmp_723_fu_18157_p3;

assign zext_ln377_95_fu_20856_p1 = tmp_729_reg_41789;

assign zext_ln377_96_fu_21005_p1 = tmp_735_reg_41818;

assign zext_ln377_97_fu_21154_p1 = tmp_741_reg_41847;

assign zext_ln377_98_fu_21303_p1 = tmp_747_reg_41876;

assign zext_ln377_99_fu_21448_p1 = tmp_753_reg_41905;

assign zext_ln377_fu_17311_p1 = tmp_fu_17303_p3;

endmodule //motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config5_s
