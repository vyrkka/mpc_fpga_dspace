module motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config8_s (
        ap_clk,
        ap_rst,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [31:0] p_read;
input  [31:0] p_read1;
input  [31:0] p_read2;
input  [31:0] p_read3;
input  [31:0] p_read4;
input  [31:0] p_read5;
input  [31:0] p_read6;
input  [31:0] p_read7;
input  [31:0] p_read8;
output  [31:0] ap_return_0;
output  [31:0] ap_return_1;
output  [31:0] ap_return_2;
output  [31:0] ap_return_3;
output  [31:0] ap_return_4;
output  [31:0] ap_return_5;
output  [31:0] ap_return_6;
output  [31:0] ap_return_7;
output  [31:0] ap_return_8;
input   ap_ce;

reg[31:0] ap_return_0;
reg[31:0] ap_return_1;
reg[31:0] ap_return_2;
reg[31:0] ap_return_3;
reg[31:0] ap_return_4;
reg[31:0] ap_return_5;
reg[31:0] ap_return_6;
reg[31:0] ap_return_7;
reg[31:0] ap_return_8;

wire   [46:0] r_V_fu_519_p2;
reg   [46:0] r_V_reg_7439;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [41:0] r_V_1_fu_470_p2;
reg   [41:0] r_V_1_reg_7443;
wire   [44:0] r_V_3_fu_510_p2;
reg   [44:0] r_V_3_reg_7447;
wire   [42:0] r_V_4_fu_526_p2;
reg   [42:0] r_V_4_reg_7451;
wire   [42:0] r_V_5_fu_500_p2;
reg   [42:0] r_V_5_reg_7455;
wire   [56:0] r_V_7_fu_537_p2;
reg   [56:0] r_V_7_reg_7459;
wire   [44:0] r_V_8_fu_514_p2;
reg   [44:0] r_V_8_reg_7463;
wire   [42:0] r_V_9_fu_503_p2;
reg   [42:0] r_V_9_reg_7467;
wire   [44:0] r_V_10_fu_548_p2;
reg   [44:0] r_V_10_reg_7471;
wire   [44:0] r_V_11_fu_478_p2;
reg   [44:0] r_V_11_reg_7475;
wire   [41:0] r_V_12_fu_489_p2;
reg   [41:0] r_V_12_reg_7479;
wire   [42:0] r_V_13_fu_501_p2;
reg   [42:0] r_V_13_reg_7483;
wire   [44:0] r_V_14_fu_546_p2;
reg   [44:0] r_V_14_reg_7487;
wire   [42:0] r_V_15_fu_482_p2;
reg   [42:0] r_V_15_reg_7491;
wire   [43:0] r_V_16_fu_492_p2;
reg   [43:0] r_V_16_reg_7495;
wire   [41:0] r_V_17_fu_485_p2;
reg   [41:0] r_V_17_reg_7499;
wire   [42:0] r_V_18_fu_481_p2;
reg   [42:0] r_V_18_reg_7503;
wire   [42:0] r_V_19_fu_473_p2;
reg   [42:0] r_V_19_reg_7507;
wire   [37:0] r_V_20_fu_515_p2;
reg   [37:0] r_V_20_reg_7511;
wire   [44:0] r_V_22_fu_535_p2;
reg   [44:0] r_V_22_reg_7515;
wire   [42:0] r_V_23_fu_518_p2;
reg   [42:0] r_V_23_reg_7519;
wire   [55:0] r_V_24_fu_508_p2;
reg   [55:0] r_V_24_reg_11671;
wire   [43:0] r_V_25_fu_497_p2;
reg   [43:0] r_V_25_reg_11675;
wire   [42:0] r_V_26_fu_490_p2;
reg   [42:0] r_V_26_reg_11679;
wire   [43:0] r_V_27_fu_541_p2;
reg   [43:0] r_V_27_reg_11683;
wire   [42:0] r_V_28_fu_521_p2;
reg   [42:0] r_V_28_reg_11687;
wire   [40:0] r_V_29_fu_538_p2;
reg   [40:0] r_V_29_reg_11691;
wire   [40:0] r_V_30_fu_488_p2;
reg   [40:0] r_V_30_reg_11695;
wire   [45:0] r_V_31_fu_496_p2;
reg   [45:0] r_V_31_reg_11699;
wire   [55:0] r_V_32_fu_499_p2;
reg   [55:0] r_V_32_reg_11703;
wire   [50:0] r_V_33_fu_527_p2;
reg   [50:0] r_V_33_reg_11707;
wire   [43:0] r_V_34_fu_509_p2;
reg   [43:0] r_V_34_reg_11711;
wire   [41:0] r_V_35_fu_476_p2;
reg   [41:0] r_V_35_reg_11715;
wire   [42:0] r_V_37_fu_494_p2;
reg   [42:0] r_V_37_reg_11719;
wire   [43:0] r_V_38_fu_498_p2;
reg   [43:0] r_V_38_reg_11723;
wire   [42:0] r_V_39_fu_505_p2;
reg   [42:0] r_V_39_reg_11727;
wire   [44:0] r_V_40_fu_512_p2;
reg   [44:0] r_V_40_reg_11731;
wire   [52:0] r_V_41_fu_472_p2;
reg   [52:0] r_V_41_reg_11735;
wire   [42:0] r_V_43_fu_531_p2;
reg   [42:0] r_V_43_reg_14203;
wire   [41:0] r_V_44_fu_520_p2;
reg   [41:0] r_V_44_reg_14207;
wire   [44:0] r_V_45_fu_506_p2;
reg   [44:0] r_V_45_reg_14211;
wire   [43:0] r_V_46_fu_530_p2;
reg   [43:0] r_V_46_reg_14215;
wire   [42:0] r_V_47_fu_471_p2;
reg   [42:0] r_V_47_reg_14219;
wire   [42:0] r_V_49_fu_480_p2;
reg   [42:0] r_V_49_reg_14223;
wire   [42:0] r_V_51_fu_491_p2;
reg   [42:0] r_V_51_reg_14227;
wire   [41:0] r_V_52_fu_523_p2;
reg   [41:0] r_V_52_reg_14231;
wire   [43:0] r_V_53_fu_534_p2;
reg   [43:0] r_V_53_reg_14235;
wire   [44:0] r_V_54_fu_493_p2;
reg   [44:0] r_V_54_reg_14239;
wire   [44:0] r_V_55_fu_540_p2;
reg   [44:0] r_V_55_reg_14243;
wire   [43:0] r_V_56_fu_549_p2;
reg   [43:0] r_V_56_reg_14247;
wire   [44:0] r_V_57_fu_504_p2;
reg   [44:0] r_V_57_reg_14251;
wire   [43:0] r_V_59_fu_532_p2;
reg   [43:0] r_V_59_reg_14255;
wire   [41:0] r_V_60_fu_474_p2;
reg   [41:0] r_V_60_reg_16179;
wire   [42:0] r_V_61_fu_543_p2;
reg   [42:0] r_V_61_reg_16183;
wire   [43:0] r_V_62_fu_477_p2;
reg   [43:0] r_V_62_reg_16187;
wire   [41:0] r_V_63_fu_545_p2;
reg   [41:0] r_V_63_reg_16191;
wire   [43:0] r_V_64_fu_533_p2;
reg   [43:0] r_V_64_reg_16195;
wire   [42:0] r_V_66_fu_511_p2;
reg   [42:0] r_V_66_reg_16199;
wire   [43:0] r_V_67_fu_522_p2;
reg   [43:0] r_V_67_reg_16203;
wire   [41:0] r_V_68_fu_544_p2;
reg   [41:0] r_V_68_reg_16207;
wire   [43:0] r_V_69_fu_529_p2;
reg   [43:0] r_V_69_reg_16211;
wire   [42:0] r_V_70_fu_516_p2;
reg   [42:0] r_V_70_reg_16215;
wire   [41:0] r_V_71_fu_517_p2;
reg   [41:0] r_V_71_reg_16219;
wire   [42:0] r_V_72_fu_525_p2;
reg   [42:0] r_V_72_reg_16223;
wire   [40:0] r_V_74_fu_495_p2;
reg   [40:0] r_V_74_reg_16227;
wire   [39:0] r_V_75_fu_539_p2;
reg   [39:0] r_V_75_reg_16231;
wire   [45:0] r_V_76_fu_484_p2;
reg   [45:0] r_V_76_reg_16235;
wire   [53:0] r_V_77_fu_486_p2;
reg   [53:0] r_V_77_reg_16239;
reg  signed [31:0] p_read_18_reg_40258;
reg  signed [31:0] p_read_18_reg_40258_pp0_iter1_reg;
reg  signed [31:0] p_read_18_reg_40258_pp0_iter2_reg;
reg  signed [31:0] p_read_19_reg_40271;
reg  signed [31:0] p_read_19_reg_40271_pp0_iter1_reg;
reg  signed [31:0] p_read_19_reg_40271_pp0_iter2_reg;
reg  signed [31:0] p_read_20_reg_40279;
reg  signed [31:0] p_read_20_reg_40279_pp0_iter1_reg;
reg  signed [31:0] p_read_21_reg_40289;
reg  signed [31:0] p_read_21_reg_40289_pp0_iter1_reg;
reg  signed [31:0] p_read_22_reg_40302;
reg  signed [31:0] p_read_23_reg_40314;
reg   [0:0] p_Result_s_reg_40323;
reg   [0:0] p_Result_1_reg_40329;
wire  signed [23:0] p_Val2_2_fu_16325_p2;
reg  signed [23:0] p_Val2_2_reg_40335;
reg   [0:0] p_Result_2_reg_40340;
reg   [0:0] Range2_all_ones_reg_40347;
reg   [0:0] p_Result_3_reg_40354;
reg   [0:0] p_Result_4_reg_40360;
wire  signed [18:0] p_Val2_5_fu_16389_p2;
reg  signed [18:0] p_Val2_5_reg_40366;
reg   [0:0] p_Result_5_reg_40371;
reg   [0:0] Range2_all_ones_1_reg_40378;
wire  signed [15:0] p_Val2_8_fu_16489_p2;
reg  signed [15:0] p_Val2_8_reg_40385;
wire   [0:0] overflow_2_fu_16591_p2;
reg   [0:0] overflow_2_reg_40390;
wire   [0:0] or_ln346_2_fu_16621_p2;
reg   [0:0] or_ln346_2_reg_40395;
reg   [0:0] p_Result_9_reg_40400;
reg   [0:0] p_Result_10_reg_40406;
wire  signed [21:0] p_Val2_11_fu_16669_p2;
reg  signed [21:0] p_Val2_11_reg_40412;
reg   [0:0] p_Result_11_reg_40417;
reg   [0:0] Range2_all_ones_3_reg_40424;
reg   [0:0] p_Result_12_reg_40431;
reg   [0:0] p_Result_13_reg_40437;
wire  signed [19:0] p_Val2_14_fu_16733_p2;
reg  signed [19:0] p_Val2_14_reg_40443;
reg   [0:0] p_Result_14_reg_40448;
reg   [0:0] Range2_all_ones_4_reg_40455;
reg   [0:0] p_Result_15_reg_40462;
reg   [0:0] p_Result_16_reg_40468;
wire  signed [19:0] p_Val2_17_fu_16797_p2;
reg  signed [19:0] p_Val2_17_reg_40474;
reg   [0:0] p_Result_17_reg_40479;
reg   [0:0] Range2_all_ones_5_reg_40486;
wire  signed [15:0] p_Val2_20_fu_16867_p2;
reg  signed [15:0] p_Val2_20_reg_40493;
wire   [0:0] overflow_6_fu_16969_p2;
reg   [0:0] overflow_6_reg_40498;
wire   [0:0] or_ln346_6_fu_16999_p2;
reg   [0:0] or_ln346_6_reg_40503;
reg   [0:0] p_Result_21_reg_40508;
reg   [0:0] p_Result_22_reg_40514;
wire   [31:0] p_Val2_23_fu_17043_p2;
reg   [31:0] p_Val2_23_reg_40520;
reg   [0:0] p_Result_23_reg_40525;
reg   [0:0] Range2_all_ones_7_reg_40532;
reg   [0:0] p_Result_24_reg_40539;
reg   [0:0] p_Result_25_reg_40545;
wire  signed [21:0] p_Val2_26_fu_17107_p2;
reg  signed [21:0] p_Val2_26_reg_40551;
reg   [0:0] p_Result_26_reg_40556;
reg   [0:0] Range2_all_ones_8_reg_40563;
reg   [0:0] p_Result_27_reg_40570;
reg   [18:0] p_Val2_28_reg_40576;
reg   [0:0] p_Result_28_reg_40581;
reg   [0:0] tmp_54_reg_40587;
reg   [0:0] Range2_all_ones_9_reg_40592;
wire  signed [17:0] p_Val2_31_fu_17231_p2;
reg  signed [17:0] p_Val2_31_reg_40599;
wire   [0:0] overflow_10_fu_17333_p2;
reg   [0:0] overflow_10_reg_40604;
wire   [0:0] or_ln346_10_fu_17363_p2;
reg   [0:0] or_ln346_10_reg_40609;
wire  signed [13:0] p_Val2_33_fu_17403_p2;
reg  signed [13:0] p_Val2_33_reg_40614;
wire   [0:0] overflow_11_fu_17477_p2;
reg   [0:0] overflow_11_reg_40619;
wire   [0:0] or_ln346_11_fu_17507_p2;
reg   [0:0] or_ln346_11_reg_40624;
reg   [0:0] p_Result_35_reg_40629;
reg   [20:0] p_Val2_35_reg_40635;
reg   [0:0] p_Result_36_reg_40640;
reg   [0:0] tmp_69_reg_40646;
reg   [0:0] Range2_all_ones_11_reg_40651;
reg   [0:0] p_Result_38_reg_40658;
reg   [20:0] p_Val2_38_reg_40664;
reg   [0:0] p_Result_39_reg_40669;
reg   [0:0] tmp_75_reg_40675;
reg   [0:0] Range2_all_ones_12_reg_40680;
wire  signed [16:0] p_Val2_41_fu_17631_p2;
reg  signed [16:0] p_Val2_41_reg_40687;
wire   [0:0] overflow_14_fu_17705_p2;
reg   [0:0] overflow_14_reg_40692;
wire   [0:0] or_ln346_14_fu_17735_p2;
reg   [0:0] or_ln346_14_reg_40697;
reg   [0:0] p_Result_43_reg_40702;
reg   [0:0] p_Result_44_reg_40708;
wire  signed [18:0] p_Val2_44_fu_17783_p2;
reg  signed [18:0] p_Val2_44_reg_40714;
reg   [0:0] p_Result_45_reg_40719;
reg   [0:0] Range2_all_ones_13_reg_40726;
reg   [0:0] p_Result_46_reg_40733;
reg   [18:0] p_Val2_46_reg_40739;
reg   [0:0] p_Result_47_reg_40744;
reg   [0:0] tmp_90_reg_40750;
reg   [0:0] Range2_all_ones_14_reg_40755;
reg   [0:0] p_Result_49_reg_40762;
reg   [20:0] p_Val2_49_reg_40768;
reg   [0:0] p_Result_50_reg_40773;
reg   [0:0] tmp_96_reg_40779;
reg   [0:0] Range2_all_ones_15_reg_40784;
reg   [0:0] p_Result_52_reg_40791;
reg   [18:0] p_Val2_52_reg_40797;
reg   [0:0] p_Result_53_reg_40802;
reg   [0:0] tmp_102_reg_40808;
reg   [0:0] Range2_all_ones_16_reg_40813;
reg   [0:0] p_Result_55_reg_40820;
reg   [19:0] p_Val2_55_reg_40826;
reg   [0:0] p_Result_56_reg_40831;
reg   [0:0] tmp_108_reg_40837;
reg   [0:0] Range2_all_ones_17_reg_40842;
reg   [0:0] p_Result_58_reg_40849;
reg   [17:0] p_Val2_58_reg_40855;
reg   [0:0] p_Result_59_reg_40860;
reg   [0:0] tmp_114_reg_40866;
reg   [0:0] Range2_all_ones_18_reg_40871;
reg   [0:0] p_Result_61_reg_40878;
reg   [18:0] p_Val2_61_reg_40884;
reg   [0:0] p_Result_62_reg_40889;
reg   [0:0] tmp_120_reg_40895;
reg   [0:0] Range2_all_ones_19_reg_40900;
reg   [0:0] p_Result_64_reg_40907;
reg   [18:0] p_Val2_64_reg_40913;
reg   [0:0] p_Result_65_reg_40918;
reg   [0:0] tmp_126_reg_40924;
reg   [0:0] Range2_all_ones_20_reg_40929;
reg   [0:0] p_Result_67_reg_40936;
reg   [13:0] p_Val2_67_reg_40942;
reg   [0:0] p_Result_68_reg_40947;
reg   [0:0] tmp_132_reg_40953;
reg   [0:0] Range2_all_ones_21_reg_40958;
wire  signed [15:0] p_Val2_71_fu_18241_p2;
reg  signed [15:0] p_Val2_71_reg_40965;
wire   [0:0] overflow_24_fu_18343_p2;
reg   [0:0] overflow_24_reg_40970;
wire   [0:0] or_ln346_24_fu_18373_p2;
reg   [0:0] or_ln346_24_reg_40975;
reg   [0:0] p_Result_73_reg_40980;
reg   [20:0] p_Val2_73_reg_40986;
reg   [0:0] p_Result_74_reg_40991;
reg   [0:0] tmp_144_reg_40997;
reg   [0:0] Range2_all_ones_23_reg_41002;
reg   [0:0] p_Result_76_reg_41009;
reg   [18:0] p_Val2_76_reg_41015;
reg   [0:0] p_Result_77_reg_41020;
reg   [0:0] tmp_150_reg_41026;
reg   [0:0] Range2_all_ones_24_reg_41031;
reg   [0:0] tmp_264_reg_41038;
reg   [0:0] tmp_264_reg_41038_pp0_iter1_reg;
wire  signed [19:0] p_Val2_53_fu_20321_p2;
reg  signed [19:0] p_Val2_53_reg_41043;
wire   [0:0] overflow_18_fu_20409_p2;
reg   [0:0] overflow_18_reg_41048;
wire   [0:0] or_ln346_18_fu_20438_p2;
reg   [0:0] or_ln346_18_reg_41053;
wire  signed [20:0] p_Val2_56_fu_20450_p2;
reg  signed [20:0] p_Val2_56_reg_41058;
wire   [0:0] overflow_19_fu_20538_p2;
reg   [0:0] overflow_19_reg_41063;
wire   [0:0] or_ln346_19_fu_20567_p2;
reg   [0:0] or_ln346_19_reg_41068;
wire  signed [19:0] p_Val2_62_fu_20728_p2;
reg  signed [19:0] p_Val2_62_reg_41073;
wire   [0:0] overflow_21_fu_20816_p2;
reg   [0:0] overflow_21_reg_41078;
wire   [0:0] or_ln346_21_fu_20845_p2;
reg   [0:0] or_ln346_21_reg_41083;
wire  signed [19:0] p_Val2_65_fu_20857_p2;
reg  signed [19:0] p_Val2_65_reg_41088;
wire   [0:0] overflow_22_fu_20945_p2;
reg   [0:0] overflow_22_reg_41093;
wire   [0:0] or_ln346_22_fu_20974_p2;
reg   [0:0] or_ln346_22_reg_41098;
wire  signed [14:0] p_Val2_68_fu_20986_p2;
reg  signed [14:0] p_Val2_68_reg_41103;
wire   [0:0] overflow_23_fu_21074_p2;
reg   [0:0] overflow_23_reg_41108;
wire   [0:0] or_ln346_23_fu_21103_p2;
reg   [0:0] or_ln346_23_reg_41113;
wire  signed [21:0] p_Val2_74_fu_21132_p2;
reg  signed [21:0] p_Val2_74_reg_41118;
wire   [0:0] overflow_25_fu_21220_p2;
reg   [0:0] overflow_25_reg_41123;
wire   [0:0] or_ln346_25_fu_21249_p2;
reg   [0:0] or_ln346_25_reg_41128;
wire  signed [19:0] p_Val2_77_fu_21261_p2;
reg  signed [19:0] p_Val2_77_reg_41133;
wire   [0:0] overflow_26_fu_21349_p2;
reg   [0:0] overflow_26_reg_41138;
wire   [0:0] or_ln346_26_fu_21378_p2;
reg   [0:0] or_ln346_26_reg_41143;
reg   [0:0] p_Result_79_reg_41148;
reg   [0:0] p_Result_80_reg_41154;
wire   [31:0] p_Val2_80_fu_21446_p2;
reg   [31:0] p_Val2_80_reg_41160;
reg   [0:0] p_Result_81_reg_41165;
reg   [0:0] Range2_all_ones_25_reg_41172;
reg   [0:0] p_Result_82_reg_41179;
reg   [0:0] p_Result_83_reg_41185;
wire  signed [20:0] p_Val2_83_fu_21510_p2;
reg  signed [20:0] p_Val2_83_reg_41191;
reg   [0:0] p_Result_84_reg_41196;
reg   [0:0] Range2_all_ones_26_reg_41203;
reg   [0:0] p_Result_85_reg_41210;
reg   [0:0] p_Result_86_reg_41216;
wire  signed [19:0] p_Val2_86_fu_21574_p2;
reg  signed [19:0] p_Val2_86_reg_41222;
reg   [0:0] p_Result_87_reg_41227;
reg   [0:0] Range2_all_ones_27_reg_41234;
reg   [0:0] p_Result_88_reg_41241;
reg   [0:0] p_Result_89_reg_41247;
wire  signed [20:0] p_Val2_89_fu_21638_p2;
reg  signed [20:0] p_Val2_89_reg_41253;
reg   [0:0] p_Result_90_reg_41258;
reg   [0:0] Range2_all_ones_28_reg_41265;
reg   [0:0] p_Result_91_reg_41272;
reg   [0:0] p_Result_92_reg_41278;
wire  signed [19:0] p_Val2_92_fu_21702_p2;
reg  signed [19:0] p_Val2_92_reg_41284;
reg   [0:0] p_Result_93_reg_41289;
reg   [0:0] Range2_all_ones_29_reg_41296;
reg   [0:0] p_Result_94_reg_41303;
reg   [0:0] p_Result_95_reg_41309;
wire  signed [17:0] p_Val2_95_fu_21766_p2;
reg  signed [17:0] p_Val2_95_reg_41315;
reg   [0:0] p_Result_96_reg_41320;
reg   [0:0] Range2_all_ones_30_reg_41327;
reg   [0:0] p_Result_97_reg_41334;
reg   [0:0] p_Result_98_reg_41340;
wire  signed [17:0] p_Val2_98_fu_21830_p2;
reg  signed [17:0] p_Val2_98_reg_41346;
reg   [0:0] p_Result_99_reg_41351;
reg   [0:0] Range2_all_ones_31_reg_41358;
reg   [0:0] p_Result_100_reg_41365;
reg   [0:0] p_Result_101_reg_41371;
wire  signed [22:0] p_Val2_101_fu_21894_p2;
reg  signed [22:0] p_Val2_101_reg_41377;
reg   [0:0] p_Result_102_reg_41382;
reg   [0:0] Range2_all_ones_32_reg_41389;
reg   [0:0] p_Result_103_reg_41396;
reg   [0:0] p_Result_104_reg_41402;
wire   [31:0] p_Val2_104_fu_21954_p2;
reg   [31:0] p_Val2_104_reg_41408;
reg   [0:0] p_Result_105_reg_41413;
reg   [0:0] Range2_all_ones_33_reg_41420;
reg   [0:0] p_Result_106_reg_41427;
reg   [26:0] p_Val2_106_reg_41433;
reg   [0:0] p_Result_107_reg_41438;
reg   [0:0] tmp_210_reg_41444;
reg   [0:0] Range2_all_ones_34_reg_41449;
reg   [0:0] p_Result_109_reg_41456;
reg   [19:0] p_Val2_109_reg_41462;
reg   [0:0] p_Result_110_reg_41467;
reg   [0:0] tmp_216_reg_41473;
reg   [0:0] Range2_all_ones_35_reg_41478;
reg   [0:0] p_Result_112_reg_41485;
reg   [17:0] p_Val2_112_reg_41491;
reg   [0:0] p_Result_113_reg_41496;
reg   [0:0] tmp_222_reg_41502;
reg   [0:0] Range2_all_ones_36_reg_41507;
wire  signed [14:0] p_Val2_116_fu_22190_p2;
reg  signed [14:0] p_Val2_116_reg_41514;
wire   [0:0] overflow_39_fu_22292_p2;
reg   [0:0] overflow_39_reg_41519;
wire   [0:0] or_ln346_39_fu_22322_p2;
reg   [0:0] or_ln346_39_reg_41524;
reg   [0:0] p_Result_118_reg_41529;
reg   [18:0] p_Val2_118_reg_41535;
reg   [0:0] p_Result_119_reg_41540;
reg   [0:0] tmp_234_reg_41546;
reg   [0:0] Range2_all_ones_38_reg_41551;
reg   [0:0] p_Result_121_reg_41558;
reg   [19:0] p_Val2_121_reg_41564;
reg   [0:0] p_Result_122_reg_41569;
reg   [0:0] tmp_240_reg_41575;
reg   [0:0] Range2_all_ones_39_reg_41580;
reg   [0:0] p_Result_124_reg_41587;
reg   [18:0] p_Val2_124_reg_41593;
reg   [0:0] p_Result_125_reg_41598;
reg   [0:0] tmp_246_reg_41604;
reg   [0:0] Range2_all_ones_40_reg_41609;
reg   [0:0] p_Result_127_reg_41616;
reg   [20:0] p_Val2_127_reg_41622;
reg   [0:0] p_Result_128_reg_41627;
reg   [0:0] tmp_252_reg_41633;
reg   [0:0] Range2_all_ones_41_reg_41638;
reg   [0:0] p_Result_130_reg_41645;
reg   [28:0] p_Val2_130_reg_41651;
reg   [0:0] p_Result_131_reg_41656;
reg   [0:0] tmp_258_reg_41662;
reg   [0:0] Range2_all_ones_42_reg_41667;
wire  signed [31:0] lhs_9_fu_23514_p3;
reg  signed [31:0] lhs_9_reg_41674;
wire  signed [31:0] lhs_10_fu_23616_p3;
reg  signed [31:0] lhs_10_reg_41680;
wire  signed [31:0] lhs_12_fu_23820_p3;
reg  signed [31:0] lhs_12_reg_41686;
wire  signed [31:0] lhs_13_fu_23922_p3;
reg  signed [31:0] lhs_13_reg_41692;
wire  signed [31:0] lhs_14_fu_24024_p3;
reg  signed [31:0] lhs_14_reg_41698;
wire  signed [31:0] lhs_16_fu_24228_p3;
reg  signed [31:0] lhs_16_reg_41704;
wire  signed [31:0] lhs_17_fu_24330_p3;
reg  signed [31:0] lhs_17_reg_41710;
reg   [0:0] p_Result_281_reg_41716;
wire   [31:0] p_Val2_281_fu_24360_p2;
reg   [31:0] p_Val2_281_reg_41723;
reg   [0:0] p_Result_282_reg_41729;
reg   [0:0] p_Result_289_reg_41736;
wire   [31:0] p_Val2_289_fu_24396_p2;
reg   [31:0] p_Val2_289_reg_41743;
reg   [0:0] p_Result_290_reg_41749;
wire  signed [14:0] p_Val2_134_fu_26926_p2;
reg  signed [14:0] p_Val2_134_reg_41756;
wire   [0:0] overflow_45_fu_27028_p2;
reg   [0:0] overflow_45_reg_41761;
wire   [0:0] or_ln346_45_fu_27058_p2;
reg   [0:0] or_ln346_45_reg_41766;
reg   [0:0] p_Result_136_reg_41771;
reg   [0:0] p_Result_137_reg_41777;
wire  signed [19:0] p_Val2_137_fu_27106_p2;
reg  signed [19:0] p_Val2_137_reg_41783;
reg   [0:0] p_Result_138_reg_41788;
reg   [0:0] Range2_all_ones_44_reg_41795;
reg   [0:0] p_Result_139_reg_41802;
reg   [0:0] p_Result_140_reg_41808;
wire  signed [18:0] p_Val2_140_fu_27170_p2;
reg  signed [18:0] p_Val2_140_reg_41814;
reg   [0:0] p_Result_141_reg_41819;
reg   [0:0] Range2_all_ones_45_reg_41826;
reg   [0:0] p_Result_142_reg_41833;
reg   [0:0] p_Result_143_reg_41839;
wire  signed [21:0] p_Val2_143_fu_27234_p2;
reg  signed [21:0] p_Val2_143_reg_41845;
reg   [0:0] p_Result_144_reg_41850;
reg   [0:0] Range2_all_ones_46_reg_41857;
reg   [0:0] p_Result_145_reg_41864;
reg   [0:0] p_Result_146_reg_41870;
wire  signed [20:0] p_Val2_146_fu_27298_p2;
reg  signed [20:0] p_Val2_146_reg_41876;
reg   [0:0] p_Result_147_reg_41881;
reg   [0:0] Range2_all_ones_47_reg_41888;
reg   [0:0] p_Result_148_reg_41895;
reg   [0:0] p_Result_149_reg_41901;
wire  signed [19:0] p_Val2_149_fu_27362_p2;
reg  signed [19:0] p_Val2_149_reg_41907;
reg   [0:0] p_Result_150_reg_41912;
reg   [0:0] Range2_all_ones_48_reg_41919;
wire  signed [18:0] p_Val2_152_fu_27460_p2;
reg  signed [18:0] p_Val2_152_reg_41926;
wire   [0:0] overflow_51_fu_27562_p2;
reg   [0:0] overflow_51_reg_41931;
wire   [0:0] or_ln346_51_fu_27592_p2;
reg   [0:0] or_ln346_51_reg_41936;
reg   [0:0] p_Result_154_reg_41941;
reg   [0:0] p_Result_155_reg_41947;
wire  signed [19:0] p_Val2_155_fu_27640_p2;
reg  signed [19:0] p_Val2_155_reg_41953;
reg   [0:0] p_Result_156_reg_41958;
reg   [0:0] Range2_all_ones_50_reg_41965;
wire  signed [18:0] p_Val2_158_fu_27721_p2;
reg  signed [18:0] p_Val2_158_reg_41972;
wire   [0:0] overflow_53_fu_27823_p2;
reg   [0:0] overflow_53_reg_41977;
wire   [0:0] or_ln346_53_fu_27853_p2;
reg   [0:0] or_ln346_53_reg_41982;
reg   [0:0] p_Result_160_reg_41987;
reg   [18:0] p_Val2_160_reg_41993;
reg   [0:0] p_Result_161_reg_41998;
reg   [0:0] tmp_318_reg_42004;
reg   [0:0] Range2_all_ones_52_reg_42009;
reg   [0:0] p_Result_163_reg_42016;
reg   [17:0] p_Val2_163_reg_42022;
reg   [0:0] p_Result_164_reg_42027;
reg   [0:0] tmp_324_reg_42033;
reg   [0:0] Range2_all_ones_53_reg_42038;
reg   [0:0] p_Result_166_reg_42045;
reg   [19:0] p_Val2_166_reg_42051;
reg   [0:0] p_Result_167_reg_42056;
reg   [0:0] tmp_330_reg_42062;
reg   [0:0] Range2_all_ones_54_reg_42067;
reg   [0:0] p_Result_169_reg_42074;
reg   [20:0] p_Val2_169_reg_42080;
reg   [0:0] p_Result_170_reg_42085;
reg   [0:0] tmp_336_reg_42091;
reg   [0:0] Range2_all_ones_55_reg_42096;
reg   [0:0] p_Result_172_reg_42103;
reg   [20:0] p_Val2_172_reg_42109;
reg   [0:0] p_Result_173_reg_42114;
reg   [0:0] tmp_342_reg_42120;
reg   [0:0] Range2_all_ones_56_reg_42125;
reg   [0:0] p_Result_175_reg_42132;
reg   [19:0] p_Val2_175_reg_42138;
reg   [0:0] p_Result_176_reg_42143;
reg   [0:0] tmp_348_reg_42149;
reg   [0:0] Range2_all_ones_57_reg_42154;
reg   [0:0] p_Result_178_reg_42161;
reg   [20:0] p_Val2_178_reg_42167;
reg   [0:0] p_Result_179_reg_42172;
reg   [0:0] tmp_354_reg_42178;
reg   [0:0] Range2_all_ones_58_reg_42183;
wire  signed [18:0] p_Val2_182_fu_28243_p2;
reg  signed [18:0] p_Val2_182_reg_42190;
wire   [0:0] overflow_61_fu_28345_p2;
reg   [0:0] overflow_61_reg_42195;
wire   [0:0] or_ln346_61_fu_28375_p2;
reg   [0:0] or_ln346_61_reg_42200;
reg   [0:0] p_Result_184_reg_42205;
reg   [19:0] p_Val2_184_reg_42211;
reg   [0:0] p_Result_185_reg_42216;
reg   [0:0] tmp_366_reg_42222;
reg   [0:0] Range2_all_ones_60_reg_42227;
reg   [0:0] p_Result_313_reg_42234;
wire   [31:0] p_Val2_313_fu_30179_p2;
reg   [31:0] p_Val2_313_reg_42241;
reg   [0:0] p_Result_314_reg_42247;
reg   [0:0] p_Result_315_reg_42254;
wire   [31:0] p_Val2_315_fu_30215_p2;
reg   [31:0] p_Val2_315_reg_42261;
reg   [0:0] p_Result_316_reg_42267;
wire  signed [31:0] lhs_38_fu_30323_p3;
reg  signed [31:0] lhs_38_reg_42274;
reg   [0:0] p_Result_319_reg_42280;
wire   [31:0] p_Val2_319_fu_30353_p2;
reg   [31:0] p_Val2_319_reg_42287;
reg   [0:0] p_Result_320_reg_42293;
reg   [0:0] p_Result_321_reg_42300;
wire   [31:0] p_Val2_321_fu_30389_p2;
reg   [31:0] p_Val2_321_reg_42307;
reg   [0:0] p_Result_322_reg_42313;
reg   [0:0] p_Result_323_reg_42320;
wire   [31:0] p_Val2_323_fu_30425_p2;
reg   [31:0] p_Val2_323_reg_42327;
reg   [0:0] p_Result_324_reg_42333;
wire  signed [31:0] lhs_42_fu_30533_p3;
reg  signed [31:0] lhs_42_reg_42340;
reg   [0:0] p_Result_327_reg_42346;
wire   [31:0] p_Val2_327_fu_30563_p2;
reg   [31:0] p_Val2_327_reg_42353;
reg   [0:0] p_Result_328_reg_42359;
reg   [0:0] p_Result_329_reg_42366;
wire   [31:0] p_Val2_329_fu_30599_p2;
reg   [31:0] p_Val2_329_reg_42373;
reg   [0:0] p_Result_330_reg_42379;
reg   [0:0] p_Result_187_reg_42386;
reg   [0:0] p_Result_188_reg_42392;
wire  signed [18:0] p_Val2_188_fu_32682_p2;
reg  signed [18:0] p_Val2_188_reg_42398;
reg   [0:0] p_Result_189_reg_42403;
reg   [0:0] Range2_all_ones_61_reg_42410;
reg   [0:0] p_Result_190_reg_42417;
reg   [0:0] p_Result_191_reg_42423;
wire  signed [19:0] p_Val2_191_fu_32746_p2;
reg  signed [19:0] p_Val2_191_reg_42429;
reg   [0:0] p_Result_192_reg_42434;
reg   [0:0] Range2_all_ones_62_reg_42441;
reg   [0:0] p_Result_193_reg_42448;
reg   [0:0] p_Result_194_reg_42454;
wire  signed [20:0] p_Val2_194_fu_32810_p2;
reg  signed [20:0] p_Val2_194_reg_42460;
reg   [0:0] p_Result_195_reg_42465;
reg   [0:0] Range2_all_ones_63_reg_42472;
reg   [0:0] p_Result_196_reg_42479;
reg   [0:0] p_Result_197_reg_42485;
wire  signed [18:0] p_Val2_197_fu_32874_p2;
reg  signed [18:0] p_Val2_197_reg_42491;
reg   [0:0] p_Result_198_reg_42496;
reg   [0:0] Range2_all_ones_64_reg_42503;
reg   [0:0] p_Result_199_reg_42510;
reg   [0:0] p_Result_200_reg_42516;
wire  signed [20:0] p_Val2_200_fu_32938_p2;
reg  signed [20:0] p_Val2_200_reg_42522;
reg   [0:0] p_Result_201_reg_42527;
reg   [0:0] Range2_all_ones_65_reg_42534;
wire  signed [15:0] p_Val2_203_fu_33019_p2;
reg  signed [15:0] p_Val2_203_reg_42541;
wire   [0:0] overflow_68_fu_33121_p2;
reg   [0:0] overflow_68_reg_42546;
wire   [0:0] or_ln346_68_fu_33151_p2;
reg   [0:0] or_ln346_68_reg_42551;
reg   [0:0] p_Result_205_reg_42556;
reg   [0:0] p_Result_206_reg_42562;
wire  signed [19:0] p_Val2_206_fu_33199_p2;
reg  signed [19:0] p_Val2_206_reg_42568;
reg   [0:0] p_Result_207_reg_42573;
reg   [0:0] Range2_all_ones_67_reg_42580;
reg   [0:0] p_Result_208_reg_42587;
reg   [0:0] p_Result_209_reg_42593;
wire  signed [20:0] p_Val2_209_fu_33263_p2;
reg  signed [20:0] p_Val2_209_reg_42599;
reg   [0:0] p_Result_210_reg_42604;
reg   [0:0] Range2_all_ones_68_reg_42611;
reg   [0:0] p_Result_211_reg_42618;
reg   [0:0] p_Result_212_reg_42624;
wire  signed [18:0] p_Val2_212_fu_33327_p2;
reg  signed [18:0] p_Val2_212_reg_42630;
reg   [0:0] p_Result_213_reg_42635;
reg   [0:0] Range2_all_ones_69_reg_42642;
reg   [0:0] p_Result_214_reg_42649;
reg   [19:0] p_Val2_214_reg_42655;
reg   [0:0] p_Result_215_reg_42660;
reg   [0:0] tmp_426_reg_42666;
reg   [0:0] Range2_all_ones_70_reg_42671;
reg   [0:0] p_Result_217_reg_42678;
reg   [18:0] p_Val2_217_reg_42684;
reg   [0:0] p_Result_218_reg_42689;
reg   [0:0] tmp_432_reg_42695;
reg   [0:0] Range2_all_ones_71_reg_42700;
reg   [0:0] p_Result_220_reg_42707;
reg   [17:0] p_Val2_220_reg_42713;
reg   [0:0] p_Result_221_reg_42718;
reg   [0:0] tmp_438_reg_42724;
reg   [0:0] Range2_all_ones_72_reg_42729;
reg   [0:0] p_Result_223_reg_42736;
reg   [18:0] p_Val2_223_reg_42742;
reg   [0:0] p_Result_224_reg_42747;
reg   [0:0] tmp_444_reg_42753;
reg   [0:0] Range2_all_ones_73_reg_42758;
wire  signed [16:0] p_Val2_227_fu_33616_p2;
reg  signed [16:0] p_Val2_227_reg_42765;
wire   [0:0] overflow_76_fu_33718_p2;
reg   [0:0] overflow_76_reg_42770;
wire   [0:0] or_ln346_76_fu_33748_p2;
reg   [0:0] or_ln346_76_reg_42775;
reg   [0:0] p_Result_229_reg_42780;
reg   [16:0] p_Val2_229_reg_42786;
reg   [0:0] p_Result_230_reg_42791;
reg   [0:0] tmp_456_reg_42797;
reg   [0:0] Range2_all_ones_75_reg_42802;
reg   [0:0] p_Result_232_reg_42809;
reg   [15:0] p_Val2_232_reg_42815;
reg   [0:0] p_Result_233_reg_42820;
reg   [0:0] tmp_462_reg_42826;
reg   [0:0] Range2_all_ones_76_reg_42831;
reg   [0:0] p_Result_235_reg_42838;
reg   [21:0] p_Val2_235_reg_42844;
reg   [0:0] p_Result_236_reg_42849;
reg   [0:0] tmp_468_reg_42855;
reg   [0:0] Range2_all_ones_77_reg_42860;
reg   [0:0] p_Result_238_reg_42867;
reg   [29:0] p_Val2_238_reg_42873;
reg   [0:0] p_Result_239_reg_42878;
reg   [0:0] tmp_474_reg_42884;
reg   [0:0] Range2_all_ones_78_reg_42889;
wire  signed [31:0] lhs_54_fu_35336_p3;
reg  signed [31:0] lhs_54_reg_42896;
wire  signed [31:0] lhs_55_fu_35438_p3;
reg  signed [31:0] lhs_55_reg_42902;
wire  signed [31:0] lhs_56_fu_35540_p3;
reg  signed [31:0] lhs_56_reg_42908;
wire  signed [31:0] lhs_57_fu_35642_p3;
reg  signed [31:0] lhs_57_reg_42914;
wire  signed [31:0] lhs_58_fu_35744_p3;
reg  signed [31:0] lhs_58_reg_42920;
wire  signed [31:0] lhs_59_fu_35846_p3;
reg  signed [31:0] lhs_59_reg_42926;
wire  signed [31:0] lhs_60_fu_35948_p3;
reg  signed [31:0] lhs_60_reg_42932;
wire  signed [31:0] lhs_61_fu_36050_p3;
reg  signed [31:0] lhs_61_reg_42938;
wire  signed [31:0] lhs_62_fu_36152_p3;
reg  signed [31:0] lhs_62_reg_42944;
wire   [9:0] r_V_1_fu_470_p1;
wire    ap_block_pp0_stage0;
wire  signed [31:0] r_V_47_fu_471_p0;
wire  signed [42:0] sext_ln70_29_fu_26867_p1;
wire   [10:0] r_V_47_fu_471_p1;
wire   [21:0] r_V_41_fu_472_p1;
wire  signed [31:0] r_V_19_fu_473_p0;
wire  signed [42:0] sext_ln70_13_fu_17909_p1;
wire   [10:0] r_V_19_fu_473_p1;
wire  signed [31:0] r_V_60_fu_474_p0;
wire  signed [41:0] sext_ln70_37_fu_32634_p1;
wire  signed [9:0] r_V_60_fu_474_p1;
wire   [9:0] r_V_35_fu_476_p1;
wire  signed [31:0] r_V_62_fu_477_p0;
wire  signed [43:0] sext_ln70_35_fu_32623_p1;
wire   [11:0] r_V_62_fu_477_p1;
wire  signed [31:0] r_V_11_fu_478_p0;
wire  signed [44:0] sext_ln70_7_fu_17134_p1;
wire  signed [12:0] r_V_11_fu_478_p1;
wire  signed [31:0] r_V_49_fu_480_p0;
wire  signed [10:0] r_V_49_fu_480_p1;
wire  signed [31:0] r_V_18_fu_481_p0;
wire  signed [10:0] r_V_18_fu_481_p1;
wire  signed [31:0] r_V_15_fu_482_p0;
wire   [10:0] r_V_15_fu_482_p1;
wire   [13:0] r_V_76_fu_484_p1;
wire   [9:0] r_V_17_fu_485_p1;
wire   [22:0] r_V_77_fu_486_p1;
wire  signed [31:0] r_V_30_fu_488_p0;
wire  signed [40:0] sext_ln70_15_fu_21388_p1;
wire  signed [8:0] r_V_30_fu_488_p1;
wire  signed [9:0] r_V_12_fu_489_p1;
wire  signed [31:0] r_V_26_fu_490_p0;
wire  signed [42:0] sext_ln70_16_fu_21393_p1;
wire   [10:0] r_V_26_fu_490_p1;
wire   [10:0] r_V_51_fu_491_p1;
wire   [11:0] r_V_16_fu_492_p1;
wire  signed [31:0] r_V_54_fu_493_p0;
wire  signed [44:0] sext_ln70_31_fu_27859_p1;
wire  signed [12:0] r_V_54_fu_493_p1;
wire  signed [31:0] r_V_37_fu_494_p0;
wire  signed [42:0] sext_ln70_21_fu_21984_p1;
wire   [10:0] r_V_37_fu_494_p1;
wire  signed [8:0] r_V_74_fu_495_p1;
wire  signed [13:0] r_V_31_fu_496_p1;
wire  signed [31:0] r_V_25_fu_497_p0;
wire  signed [43:0] sext_ln70_17_fu_21398_p1;
wire  signed [11:0] r_V_25_fu_497_p1;
wire  signed [31:0] r_V_38_fu_498_p0;
wire  signed [43:0] sext_ln70_24_fu_21996_p1;
wire  signed [11:0] r_V_38_fu_498_p1;
wire  signed [31:0] r_V_32_fu_499_p0;
wire  signed [55:0] sext_ln70_18_fu_21403_p1;
wire  signed [24:0] r_V_32_fu_499_p1;
wire  signed [31:0] r_V_5_fu_500_p0;
wire  signed [42:0] sext_ln70_1_fu_16257_p1;
wire  signed [10:0] r_V_5_fu_500_p1;
wire  signed [31:0] r_V_13_fu_501_p0;
wire  signed [42:0] sext_ln70_8_fu_17141_p1;
wire  signed [10:0] r_V_13_fu_501_p1;
wire  signed [31:0] r_V_9_fu_503_p0;
wire   [10:0] r_V_9_fu_503_p1;
wire  signed [31:0] r_V_57_fu_504_p0;
wire  signed [12:0] r_V_57_fu_504_p1;
wire  signed [31:0] r_V_39_fu_505_p0;
wire  signed [10:0] r_V_39_fu_505_p1;
wire   [12:0] r_V_45_fu_506_p1;
wire  signed [31:0] r_V_24_fu_508_p0;
wire   [24:0] r_V_24_fu_508_p1;
wire  signed [31:0] r_V_34_fu_509_p0;
wire  signed [11:0] r_V_34_fu_509_p1;
wire  signed [31:0] r_V_3_fu_510_p0;
wire  signed [44:0] sext_ln70_2_fu_16263_p1;
wire  signed [12:0] r_V_3_fu_510_p1;
wire  signed [31:0] r_V_66_fu_511_p0;
wire  signed [42:0] sext_ln70_36_fu_32629_p1;
wire  signed [10:0] r_V_66_fu_511_p1;
wire   [12:0] r_V_40_fu_512_p1;
wire  signed [31:0] r_V_8_fu_514_p0;
wire   [12:0] r_V_8_fu_514_p1;
wire  signed [5:0] r_V_20_fu_515_p1;
wire  signed [31:0] r_V_70_fu_516_p0;
wire  signed [42:0] sext_ln70_43_fu_33369_p1;
wire   [10:0] r_V_70_fu_516_p1;
wire  signed [9:0] r_V_71_fu_517_p1;
wire  signed [31:0] r_V_23_fu_518_p0;
wire  signed [10:0] r_V_23_fu_518_p1;
wire  signed [14:0] r_V_fu_519_p1;
wire  signed [9:0] r_V_44_fu_520_p1;
wire  signed [31:0] r_V_28_fu_521_p0;
wire   [10:0] r_V_28_fu_521_p1;
wire  signed [31:0] r_V_67_fu_522_p0;
wire  signed [11:0] r_V_67_fu_522_p1;
wire  signed [9:0] r_V_52_fu_523_p1;
wire  signed [31:0] r_V_72_fu_525_p0;
wire  signed [10:0] r_V_72_fu_525_p1;
wire  signed [31:0] r_V_4_fu_526_p0;
wire  signed [10:0] r_V_4_fu_526_p1;
wire  signed [19:0] r_V_33_fu_527_p1;
wire  signed [11:0] r_V_69_fu_529_p1;
wire  signed [11:0] r_V_46_fu_530_p1;
wire  signed [31:0] r_V_43_fu_531_p0;
wire  signed [10:0] r_V_43_fu_531_p1;
wire  signed [31:0] r_V_59_fu_532_p0;
wire  signed [43:0] sext_ln70_32_fu_27865_p1;
wire  signed [11:0] r_V_59_fu_532_p1;
wire  signed [31:0] r_V_64_fu_533_p0;
wire   [11:0] r_V_64_fu_533_p1;
wire  signed [31:0] r_V_53_fu_534_p0;
wire   [11:0] r_V_53_fu_534_p1;
wire  signed [12:0] r_V_22_fu_535_p1;
wire  signed [25:0] r_V_7_fu_537_p1;
wire  signed [31:0] r_V_29_fu_538_p0;
wire  signed [8:0] r_V_29_fu_538_p1;
wire   [7:0] r_V_75_fu_539_p1;
wire  signed [31:0] r_V_55_fu_540_p0;
wire   [12:0] r_V_55_fu_540_p1;
wire  signed [31:0] r_V_27_fu_541_p0;
wire  signed [11:0] r_V_27_fu_541_p1;
wire  signed [31:0] r_V_61_fu_543_p0;
wire   [10:0] r_V_61_fu_543_p1;
wire  signed [31:0] r_V_68_fu_544_p0;
wire  signed [9:0] r_V_68_fu_544_p1;
wire  signed [31:0] r_V_63_fu_545_p0;
wire  signed [9:0] r_V_63_fu_545_p1;
wire  signed [31:0] r_V_14_fu_546_p0;
wire   [12:0] r_V_14_fu_546_p1;
wire  signed [31:0] r_V_10_fu_548_p0;
wire   [12:0] r_V_10_fu_548_p1;
wire  signed [31:0] r_V_56_fu_549_p0;
wire  signed [11:0] r_V_56_fu_549_p1;
wire  signed [31:0] trunc_ln33_fu_16244_p0;
wire  signed [31:0] trunc_ln33_1_fu_16248_p0;
wire  signed [31:0] sext_ln70_1_fu_16257_p0;
wire  signed [31:0] sext_ln70_2_fu_16263_p0;
wire  signed [31:0] sext_ln70_3_fu_16269_p0;
wire   [22:0] p_Val2_1_fu_16291_p4;
wire   [0:0] tmp_fu_16313_p3;
wire   [23:0] zext_ln377_fu_16321_p1;
wire  signed [23:0] sext_ln823_3_fu_16301_p1;
wire   [17:0] p_Val2_4_fu_16355_p4;
wire   [0:0] tmp_6_fu_16377_p3;
wire   [18:0] zext_ln377_1_fu_16385_p1;
wire  signed [18:0] sext_ln823_4_fu_16365_p1;
wire  signed [31:0] shl_ln_fu_16411_p1;
wire   [37:0] shl_ln_fu_16411_p3;
wire  signed [31:0] trunc_ln1273_fu_16423_p0;
wire   [17:0] trunc_ln1273_fu_16423_p1;
wire  signed [38:0] sext_ln70_3_fu_16269_p1;
wire  signed [38:0] sext_ln1273_fu_16419_p1;
wire   [38:0] r_V_2_fu_16435_p2;
wire   [14:0] p_Val2_7_fu_16449_p4;
wire   [23:0] trunc_ln33_1_fu_16248_p1;
wire   [23:0] trunc_ln1_fu_16427_p3;
wire   [23:0] sub_ln823_fu_16463_p2;
wire   [0:0] tmp_12_fu_16477_p3;
wire   [15:0] zext_ln377_2_fu_16485_p1;
wire  signed [15:0] sext_ln823_5_fu_16459_p1;
wire   [0:0] p_Result_8_fu_16495_p3;
wire   [0:0] p_Result_7_fu_16469_p3;
wire   [0:0] xor_ln896_4_fu_16503_p2;
wire   [0:0] xor_ln888_7_fu_16523_p2;
wire   [0:0] Range2_all_ones_2_fu_16515_p3;
wire   [0:0] or_ln888_5_fu_16529_p2;
wire   [0:0] tmp_15_fu_16541_p3;
wire   [0:0] xor_ln890_2_fu_16549_p2;
wire   [0:0] or_ln890_5_fu_16555_p2;
wire   [0:0] carry_5_fu_16509_p2;
wire   [0:0] deleted_zeros_2_fu_16535_p2;
wire   [0:0] xor_ln895_4_fu_16573_p2;
wire   [0:0] p_Result_6_fu_16441_p3;
wire   [0:0] or_ln895_2_fu_16579_p2;
wire   [0:0] xor_ln895_5_fu_16585_p2;
wire   [0:0] deleted_ones_2_fu_16561_p2;
wire   [0:0] xor_ln896_5_fu_16597_p2;
wire   [0:0] and_ln891_2_fu_16567_p2;
wire   [0:0] or_ln896_2_fu_16603_p2;
wire   [0:0] xor_ln896_245_fu_16609_p2;
wire   [0:0] underflow_2_fu_16615_p2;
wire   [20:0] p_Val2_10_fu_16635_p4;
wire   [0:0] tmp_18_fu_16657_p3;
wire   [21:0] zext_ln377_3_fu_16665_p1;
wire  signed [21:0] sext_ln823_6_fu_16645_p1;
wire   [18:0] p_Val2_13_fu_16699_p4;
wire   [0:0] tmp_24_fu_16721_p3;
wire   [19:0] zext_ln377_4_fu_16729_p1;
wire  signed [19:0] sext_ln823_7_fu_16709_p1;
wire   [18:0] p_Val2_16_fu_16763_p4;
wire   [0:0] tmp_30_fu_16785_p3;
wire   [19:0] zext_ln377_5_fu_16793_p1;
wire  signed [19:0] sext_ln823_8_fu_16773_p1;
wire   [38:0] r_V_6_fu_16819_p2;
wire   [14:0] p_Val2_19_fu_16833_p4;
wire   [0:0] tmp_36_fu_16855_p3;
wire   [15:0] zext_ln377_6_fu_16863_p1;
wire  signed [15:0] sext_ln823_9_fu_16843_p1;
wire   [0:0] p_Result_20_fu_16873_p3;
wire   [0:0] p_Result_19_fu_16847_p3;
wire   [0:0] xor_ln896_12_fu_16881_p2;
wire   [0:0] xor_ln888_15_fu_16901_p2;
wire   [0:0] Range2_all_ones_6_fu_16893_p3;
wire   [0:0] or_ln888_9_fu_16907_p2;
wire   [0:0] tmp_39_fu_16919_p3;
wire   [0:0] xor_ln890_6_fu_16927_p2;
wire   [0:0] or_ln890_9_fu_16933_p2;
wire   [0:0] carry_13_fu_16887_p2;
wire   [0:0] deleted_zeros_6_fu_16913_p2;
wire   [0:0] xor_ln895_12_fu_16951_p2;
wire   [0:0] p_Result_18_fu_16825_p3;
wire   [0:0] or_ln895_6_fu_16957_p2;
wire   [0:0] xor_ln895_13_fu_16963_p2;
wire   [0:0] deleted_ones_6_fu_16939_p2;
wire   [0:0] xor_ln896_13_fu_16975_p2;
wire   [0:0] and_ln891_6_fu_16945_p2;
wire   [0:0] or_ln896_6_fu_16981_p2;
wire   [0:0] xor_ln896_249_fu_16987_p2;
wire   [0:0] underflow_6_fu_16993_p2;
wire   [0:0] tmp_42_fu_17031_p3;
wire   [31:0] zext_ln377_7_fu_17039_p1;
wire   [31:0] p_Val2_22_fu_17013_p4;
wire   [20:0] p_Val2_25_fu_17073_p4;
wire   [0:0] tmp_48_fu_17095_p3;
wire   [21:0] zext_ln377_8_fu_17103_p1;
wire  signed [21:0] sext_ln823_10_fu_17083_p1;
wire  signed [31:0] sext_ln70_7_fu_17134_p0;
wire  signed [31:0] sext_ln70_8_fu_17141_p0;
wire  signed [31:0] p_Result_30_fu_17189_p1;
wire  signed [31:0] p_Val2_30_fu_17197_p1;
wire   [16:0] p_Val2_30_fu_17197_p4;
wire  signed [31:0] p_Result_31_fu_17211_p1;
wire  signed [31:0] tmp_60_fu_17219_p1;
wire   [0:0] tmp_60_fu_17219_p3;
wire   [17:0] zext_ln377_10_fu_17227_p1;
wire  signed [17:0] sext_ln823_fu_17207_p1;
wire   [0:0] p_Result_32_fu_17237_p3;
wire  signed [31:0] Range2_all_ones_10_fu_17251_p1;
wire   [0:0] p_Result_31_fu_17211_p3;
wire   [0:0] xor_ln888_fu_17259_p2;
wire  signed [31:0] tmp_63_fu_17271_p1;
wire   [0:0] tmp_63_fu_17271_p3;
wire   [0:0] or_ln888_fu_17265_p2;
wire   [0:0] xor_ln890_10_fu_17279_p2;
wire   [0:0] Range2_all_ones_10_fu_17251_p3;
wire   [0:0] or_ln890_fu_17285_p2;
wire   [0:0] xor_ln896_20_fu_17245_p2;
wire   [0:0] and_ln891_81_fu_17297_p2;
wire   [0:0] xor_ln895_23_fu_17309_p2;
wire   [0:0] xor_ln895_20_fu_17315_p2;
wire   [0:0] p_Result_30_fu_17189_p3;
wire   [0:0] or_ln895_10_fu_17321_p2;
wire   [0:0] xor_ln895_21_fu_17327_p2;
wire   [0:0] deleted_ones_10_fu_17291_p2;
wire   [0:0] xor_ln896_21_fu_17339_p2;
wire   [0:0] and_ln891_10_fu_17303_p2;
wire   [0:0] or_ln896_10_fu_17345_p2;
wire   [0:0] xor_ln896_253_fu_17351_p2;
wire   [0:0] underflow_10_fu_17357_p2;
wire  signed [31:0] p_Val2_32_fu_17369_p1;
wire   [12:0] p_Val2_32_fu_17369_p4;
wire  signed [31:0] p_Result_33_fu_17383_p1;
wire  signed [31:0] tmp_65_fu_17391_p1;
wire   [0:0] tmp_65_fu_17391_p3;
wire   [13:0] zext_ln377_11_fu_17399_p1;
wire  signed [13:0] sext_ln823_1_fu_17379_p1;
wire   [0:0] p_Result_34_fu_17409_p3;
wire   [0:0] p_Result_33_fu_17383_p3;
wire   [0:0] xor_ln888_2_fu_17423_p2;
wire   [0:0] or_ln888_1_fu_17429_p2;
wire   [0:0] or_ln890_1_fu_17435_p2;
wire   [0:0] xor_ln896_22_fu_17417_p2;
wire   [0:0] and_ln891_82_fu_17447_p2;
wire   [0:0] xor_ln895_29_fu_17459_p2;
wire   [0:0] xor_ln895_22_fu_17465_p2;
wire   [0:0] or_ln895_11_fu_17471_p2;
wire   [0:0] deleted_ones_11_fu_17441_p2;
wire   [0:0] xor_ln896_23_fu_17483_p2;
wire   [0:0] and_ln891_11_fu_17453_p2;
wire   [0:0] or_ln896_11_fu_17489_p2;
wire   [0:0] xor_ln896_254_fu_17495_p2;
wire   [0:0] underflow_11_fu_17501_p2;
wire  signed [31:0] p_Val2_40_fu_17597_p1;
wire   [15:0] p_Val2_40_fu_17597_p4;
wire  signed [31:0] p_Result_41_fu_17611_p1;
wire  signed [31:0] tmp_80_fu_17619_p1;
wire   [0:0] tmp_80_fu_17619_p3;
wire   [16:0] zext_ln377_14_fu_17627_p1;
wire  signed [16:0] sext_ln823_2_fu_17607_p1;
wire   [0:0] p_Result_42_fu_17637_p3;
wire   [0:0] p_Result_41_fu_17611_p3;
wire   [0:0] xor_ln888_4_fu_17651_p2;
wire   [0:0] or_ln888_2_fu_17657_p2;
wire   [0:0] or_ln890_2_fu_17663_p2;
wire   [0:0] xor_ln896_28_fu_17645_p2;
wire   [0:0] and_ln891_83_fu_17675_p2;
wire   [0:0] xor_ln895_243_fu_17687_p2;
wire   [0:0] xor_ln895_28_fu_17693_p2;
wire   [0:0] or_ln895_14_fu_17699_p2;
wire   [0:0] deleted_ones_14_fu_17669_p2;
wire   [0:0] xor_ln896_29_fu_17711_p2;
wire   [0:0] and_ln891_14_fu_17681_p2;
wire   [0:0] or_ln896_14_fu_17717_p2;
wire   [0:0] xor_ln896_257_fu_17723_p2;
wire   [0:0] underflow_14_fu_17729_p2;
wire   [17:0] p_Val2_43_fu_17749_p4;
wire   [0:0] tmp_84_fu_17771_p3;
wire   [18:0] zext_ln377_15_fu_17779_p1;
wire  signed [18:0] sext_ln823_14_fu_17759_p1;
wire  signed [31:0] sext_ln70_13_fu_17909_p0;
wire  signed [31:0] shl_ln1273_1_fu_18169_p1;
wire   [37:0] shl_ln1273_1_fu_18169_p3;
wire  signed [31:0] shl_ln1273_2_fu_18181_p1;
wire   [33:0] shl_ln1273_2_fu_18181_p3;
wire  signed [38:0] sext_ln1273_1_fu_18177_p1;
wire  signed [38:0] sext_ln1273_2_fu_18189_p1;
wire   [38:0] r_V_21_fu_18193_p2;
wire   [14:0] p_Val2_70_fu_18207_p4;
wire   [0:0] tmp_138_fu_18229_p3;
wire   [15:0] zext_ln377_24_fu_18237_p1;
wire  signed [15:0] sext_ln823_23_fu_18217_p1;
wire   [0:0] p_Result_72_fu_18247_p3;
wire   [0:0] p_Result_71_fu_18221_p3;
wire   [0:0] xor_ln896_48_fu_18255_p2;
wire   [0:0] xor_ln888_45_fu_18275_p2;
wire   [0:0] Range2_all_ones_22_fu_18267_p3;
wire   [0:0] or_ln888_24_fu_18281_p2;
wire   [0:0] tmp_141_fu_18293_p3;
wire   [0:0] xor_ln890_22_fu_18301_p2;
wire   [0:0] or_ln890_24_fu_18307_p2;
wire   [0:0] carry_46_fu_18261_p2;
wire   [0:0] deleted_zeros_21_fu_18287_p2;
wire   [0:0] xor_ln895_48_fu_18325_p2;
wire   [0:0] p_Result_70_fu_18199_p3;
wire   [0:0] or_ln895_24_fu_18331_p2;
wire   [0:0] xor_ln895_49_fu_18337_p2;
wire   [0:0] deleted_ones_24_fu_18313_p2;
wire   [0:0] xor_ln896_49_fu_18349_p2;
wire   [0:0] and_ln891_24_fu_18319_p2;
wire   [0:0] or_ln896_24_fu_18355_p2;
wire   [0:0] xor_ln896_267_fu_18361_p2;
wire   [0:0] underflow_24_fu_18367_p2;
wire  signed [31:0] trunc_ln1273_2_fu_18463_p0;
wire   [18:0] trunc_ln1273_2_fu_18463_p1;
wire   [23:0] trunc_ln33_fu_16244_p1;
wire   [23:0] trunc_ln1273_1_fu_18467_p3;
wire   [23:0] sub_ln823_1_fu_18475_p2;
wire   [0:0] xor_ln896_fu_18492_p2;
wire   [0:0] xor_ln888_1_fu_18502_p2;
wire   [0:0] or_ln888_3_fu_18507_p2;
wire   [0:0] tmp_3_fu_18517_p3;
wire   [0:0] xor_ln890_fu_18525_p2;
wire   [0:0] or_ln890_3_fu_18531_p2;
wire   [0:0] carry_1_fu_18497_p2;
wire   [0:0] deleted_zeros_fu_18512_p2;
wire   [0:0] xor_ln895_fu_18547_p2;
wire   [0:0] or_ln895_fu_18553_p2;
wire   [0:0] xor_ln895_1_fu_18558_p2;
wire   [0:0] deleted_ones_fu_18537_p2;
wire   [0:0] xor_ln896_1_fu_18569_p2;
wire   [0:0] and_ln891_fu_18542_p2;
wire   [0:0] or_ln896_fu_18575_p2;
wire   [0:0] xor_ln896_243_fu_18581_p2;
wire   [0:0] overflow_fu_18563_p2;
wire   [0:0] underflow_fu_18587_p2;
wire   [0:0] or_ln346_fu_18600_p2;
wire   [31:0] select_ln346_fu_18592_p3;
wire  signed [31:0] sext_ln856_3_fu_18489_p1;
wire   [0:0] xor_ln896_2_fu_18617_p2;
wire   [0:0] xor_ln888_5_fu_18627_p2;
wire   [0:0] or_ln888_4_fu_18632_p2;
wire   [0:0] tmp_9_fu_18642_p3;
wire   [0:0] xor_ln890_1_fu_18650_p2;
wire   [0:0] or_ln890_4_fu_18656_p2;
wire   [0:0] carry_3_fu_18622_p2;
wire   [0:0] deleted_zeros_1_fu_18637_p2;
wire   [0:0] xor_ln895_2_fu_18672_p2;
wire   [0:0] or_ln895_1_fu_18678_p2;
wire   [0:0] xor_ln895_3_fu_18683_p2;
wire   [0:0] deleted_ones_1_fu_18662_p2;
wire   [0:0] xor_ln896_3_fu_18694_p2;
wire   [0:0] and_ln891_1_fu_18667_p2;
wire   [0:0] or_ln896_1_fu_18700_p2;
wire   [0:0] xor_ln896_244_fu_18706_p2;
wire   [0:0] overflow_1_fu_18688_p2;
wire   [0:0] underflow_1_fu_18712_p2;
wire   [0:0] or_ln346_1_fu_18725_p2;
wire   [31:0] select_ln346_2_fu_18717_p3;
wire  signed [31:0] sext_ln856_4_fu_18614_p1;
wire   [31:0] select_ln346_4_fu_18742_p3;
wire  signed [31:0] sext_ln856_5_fu_18739_p1;
wire   [0:0] xor_ln896_6_fu_18759_p2;
wire   [0:0] xor_ln888_9_fu_18769_p2;
wire   [0:0] or_ln888_6_fu_18774_p2;
wire   [0:0] tmp_21_fu_18784_p3;
wire   [0:0] xor_ln890_3_fu_18792_p2;
wire   [0:0] or_ln890_6_fu_18798_p2;
wire   [0:0] carry_7_fu_18764_p2;
wire   [0:0] deleted_zeros_3_fu_18779_p2;
wire   [0:0] xor_ln895_6_fu_18814_p2;
wire   [0:0] or_ln895_3_fu_18820_p2;
wire   [0:0] xor_ln895_7_fu_18825_p2;
wire   [0:0] deleted_ones_3_fu_18804_p2;
wire   [0:0] xor_ln896_7_fu_18836_p2;
wire   [0:0] and_ln891_3_fu_18809_p2;
wire   [0:0] or_ln896_3_fu_18842_p2;
wire   [0:0] xor_ln896_246_fu_18848_p2;
wire   [0:0] overflow_3_fu_18830_p2;
wire   [0:0] underflow_3_fu_18854_p2;
wire   [0:0] or_ln346_3_fu_18867_p2;
wire   [31:0] select_ln346_6_fu_18859_p3;
wire  signed [31:0] sext_ln856_6_fu_18756_p1;
wire   [0:0] xor_ln896_8_fu_18884_p2;
wire   [0:0] xor_ln888_11_fu_18894_p2;
wire   [0:0] or_ln888_7_fu_18899_p2;
wire   [0:0] tmp_27_fu_18909_p3;
wire   [0:0] xor_ln890_4_fu_18917_p2;
wire   [0:0] or_ln890_7_fu_18923_p2;
wire   [0:0] carry_9_fu_18889_p2;
wire   [0:0] deleted_zeros_4_fu_18904_p2;
wire   [0:0] xor_ln895_8_fu_18939_p2;
wire   [0:0] or_ln895_4_fu_18945_p2;
wire   [0:0] xor_ln895_9_fu_18950_p2;
wire   [0:0] deleted_ones_4_fu_18929_p2;
wire   [0:0] xor_ln896_9_fu_18961_p2;
wire   [0:0] and_ln891_4_fu_18934_p2;
wire   [0:0] or_ln896_4_fu_18967_p2;
wire   [0:0] xor_ln896_247_fu_18973_p2;
wire   [0:0] overflow_4_fu_18955_p2;
wire   [0:0] underflow_4_fu_18979_p2;
wire   [0:0] or_ln346_4_fu_18992_p2;
wire   [31:0] select_ln346_8_fu_18984_p3;
wire  signed [31:0] sext_ln856_7_fu_18881_p1;
wire   [0:0] xor_ln896_10_fu_19009_p2;
wire   [0:0] xor_ln888_13_fu_19019_p2;
wire   [0:0] or_ln888_8_fu_19024_p2;
wire   [0:0] tmp_33_fu_19034_p3;
wire   [0:0] xor_ln890_5_fu_19042_p2;
wire   [0:0] or_ln890_8_fu_19048_p2;
wire   [0:0] carry_11_fu_19014_p2;
wire   [0:0] deleted_zeros_5_fu_19029_p2;
wire   [0:0] xor_ln895_10_fu_19064_p2;
wire   [0:0] or_ln895_5_fu_19070_p2;
wire   [0:0] xor_ln895_11_fu_19075_p2;
wire   [0:0] deleted_ones_5_fu_19054_p2;
wire   [0:0] xor_ln896_11_fu_19086_p2;
wire   [0:0] and_ln891_5_fu_19059_p2;
wire   [0:0] or_ln896_5_fu_19092_p2;
wire   [0:0] xor_ln896_248_fu_19098_p2;
wire   [0:0] overflow_5_fu_19080_p2;
wire   [0:0] underflow_5_fu_19104_p2;
wire   [0:0] or_ln346_5_fu_19117_p2;
wire   [31:0] select_ln346_10_fu_19109_p3;
wire  signed [31:0] sext_ln856_8_fu_19006_p1;
wire   [31:0] select_ln346_12_fu_19134_p3;
wire  signed [31:0] sext_ln856_9_fu_19131_p1;
wire   [0:0] xor_ln896_14_fu_19148_p2;
wire   [0:0] xor_ln888_17_fu_19158_p2;
wire   [0:0] or_ln888_10_fu_19163_p2;
wire   [0:0] tmp_45_fu_19173_p3;
wire   [0:0] xor_ln890_7_fu_19181_p2;
wire   [0:0] or_ln890_10_fu_19187_p2;
wire   [0:0] carry_15_fu_19153_p2;
wire   [0:0] deleted_zeros_7_fu_19168_p2;
wire   [0:0] xor_ln895_14_fu_19203_p2;
wire   [0:0] or_ln895_7_fu_19209_p2;
wire   [0:0] xor_ln895_15_fu_19214_p2;
wire   [0:0] deleted_ones_7_fu_19193_p2;
wire   [0:0] xor_ln896_15_fu_19225_p2;
wire   [0:0] and_ln891_7_fu_19198_p2;
wire   [0:0] or_ln896_7_fu_19231_p2;
wire   [0:0] xor_ln896_250_fu_19237_p2;
wire   [0:0] overflow_7_fu_19219_p2;
wire   [0:0] underflow_7_fu_19243_p2;
wire   [0:0] or_ln346_7_fu_19256_p2;
wire   [31:0] select_ln346_14_fu_19248_p3;
wire   [0:0] xor_ln896_16_fu_19272_p2;
wire   [0:0] xor_ln888_19_fu_19282_p2;
wire   [0:0] or_ln888_11_fu_19287_p2;
wire   [0:0] tmp_51_fu_19297_p3;
wire   [0:0] xor_ln890_8_fu_19305_p2;
wire   [0:0] or_ln890_11_fu_19311_p2;
wire   [0:0] carry_17_fu_19277_p2;
wire   [0:0] deleted_zeros_8_fu_19292_p2;
wire   [0:0] xor_ln895_16_fu_19327_p2;
wire   [0:0] or_ln895_8_fu_19333_p2;
wire   [0:0] xor_ln895_17_fu_19338_p2;
wire   [0:0] deleted_ones_8_fu_19317_p2;
wire   [0:0] xor_ln896_17_fu_19349_p2;
wire   [0:0] and_ln891_8_fu_19322_p2;
wire   [0:0] or_ln896_8_fu_19355_p2;
wire   [0:0] xor_ln896_251_fu_19361_p2;
wire   [0:0] overflow_8_fu_19343_p2;
wire   [0:0] underflow_8_fu_19367_p2;
wire   [0:0] or_ln346_8_fu_19380_p2;
wire   [31:0] select_ln346_16_fu_19372_p3;
wire  signed [31:0] sext_ln856_10_fu_19269_p1;
wire   [19:0] zext_ln377_9_fu_19397_p1;
wire  signed [19:0] sext_ln823_11_fu_19394_p1;
wire  signed [19:0] p_Val2_29_fu_19400_p2;
wire   [0:0] p_Result_29_fu_19410_p3;
wire   [0:0] xor_ln896_18_fu_19418_p2;
wire   [0:0] xor_ln888_21_fu_19429_p2;
wire   [0:0] or_ln888_12_fu_19434_p2;
wire   [0:0] tmp_57_fu_19445_p3;
wire   [0:0] xor_ln890_9_fu_19453_p2;
wire   [0:0] or_ln890_12_fu_19459_p2;
wire   [0:0] carry_19_fu_19424_p2;
wire   [0:0] deleted_zeros_9_fu_19440_p2;
wire   [0:0] xor_ln895_18_fu_19475_p2;
wire   [0:0] or_ln895_9_fu_19481_p2;
wire   [0:0] xor_ln895_19_fu_19487_p2;
wire   [0:0] deleted_ones_9_fu_19465_p2;
wire   [0:0] xor_ln896_19_fu_19498_p2;
wire   [0:0] and_ln891_9_fu_19470_p2;
wire   [0:0] or_ln896_9_fu_19504_p2;
wire   [0:0] xor_ln896_252_fu_19510_p2;
wire   [0:0] overflow_9_fu_19492_p2;
wire   [0:0] underflow_9_fu_19516_p2;
wire   [0:0] or_ln346_9_fu_19529_p2;
wire   [31:0] select_ln346_18_fu_19521_p3;
wire  signed [31:0] sext_ln856_11_fu_19406_p1;
wire   [31:0] select_ln346_20_fu_19546_p3;
wire  signed [31:0] sext_ln856_fu_19543_p1;
wire   [31:0] select_ln346_22_fu_19563_p3;
wire  signed [31:0] sext_ln856_1_fu_19560_p1;
wire   [21:0] zext_ln377_12_fu_19580_p1;
wire  signed [21:0] sext_ln823_12_fu_19577_p1;
wire  signed [21:0] p_Val2_36_fu_19583_p2;
wire   [0:0] p_Result_37_fu_19593_p3;
wire   [0:0] xor_ln896_24_fu_19601_p2;
wire   [0:0] xor_ln888_23_fu_19612_p2;
wire   [0:0] or_ln888_13_fu_19617_p2;
wire   [0:0] tmp_72_fu_19628_p3;
wire   [0:0] xor_ln890_11_fu_19636_p2;
wire   [0:0] or_ln890_13_fu_19642_p2;
wire   [0:0] carry_23_fu_19607_p2;
wire   [0:0] deleted_zeros_10_fu_19623_p2;
wire   [0:0] xor_ln895_24_fu_19658_p2;
wire   [0:0] or_ln895_12_fu_19664_p2;
wire   [0:0] xor_ln895_25_fu_19670_p2;
wire   [0:0] deleted_ones_12_fu_19648_p2;
wire   [0:0] xor_ln896_25_fu_19681_p2;
wire   [0:0] and_ln891_12_fu_19653_p2;
wire   [0:0] or_ln896_12_fu_19687_p2;
wire   [0:0] xor_ln896_255_fu_19693_p2;
wire   [0:0] overflow_12_fu_19675_p2;
wire   [0:0] underflow_12_fu_19699_p2;
wire   [0:0] or_ln346_12_fu_19712_p2;
wire   [31:0] select_ln346_24_fu_19704_p3;
wire  signed [31:0] sext_ln856_12_fu_19589_p1;
wire   [21:0] zext_ln377_13_fu_19729_p1;
wire  signed [21:0] sext_ln823_13_fu_19726_p1;
wire  signed [21:0] p_Val2_39_fu_19732_p2;
wire   [0:0] p_Result_40_fu_19742_p3;
wire   [0:0] xor_ln896_26_fu_19750_p2;
wire   [0:0] xor_ln888_25_fu_19761_p2;
wire   [0:0] or_ln888_14_fu_19766_p2;
wire   [0:0] tmp_78_fu_19777_p3;
wire   [0:0] xor_ln890_12_fu_19785_p2;
wire   [0:0] or_ln890_14_fu_19791_p2;
wire   [0:0] carry_25_fu_19756_p2;
wire   [0:0] deleted_zeros_11_fu_19772_p2;
wire   [0:0] xor_ln895_26_fu_19807_p2;
wire   [0:0] or_ln895_13_fu_19813_p2;
wire   [0:0] xor_ln895_27_fu_19819_p2;
wire   [0:0] deleted_ones_13_fu_19797_p2;
wire   [0:0] xor_ln896_27_fu_19830_p2;
wire   [0:0] and_ln891_13_fu_19802_p2;
wire   [0:0] or_ln896_13_fu_19836_p2;
wire   [0:0] xor_ln896_256_fu_19842_p2;
wire   [0:0] overflow_13_fu_19824_p2;
wire   [0:0] underflow_13_fu_19848_p2;
wire   [0:0] or_ln346_13_fu_19861_p2;
wire   [31:0] select_ln346_26_fu_19853_p3;
wire  signed [31:0] sext_ln856_13_fu_19738_p1;
wire   [31:0] select_ln346_28_fu_19878_p3;
wire  signed [31:0] sext_ln856_2_fu_19875_p1;
wire   [0:0] xor_ln896_30_fu_19895_p2;
wire   [0:0] xor_ln888_27_fu_19905_p2;
wire   [0:0] or_ln888_15_fu_19910_p2;
wire   [0:0] tmp_87_fu_19920_p3;
wire   [0:0] xor_ln890_13_fu_19928_p2;
wire   [0:0] or_ln890_15_fu_19934_p2;
wire   [0:0] carry_28_fu_19900_p2;
wire   [0:0] deleted_zeros_12_fu_19915_p2;
wire   [0:0] xor_ln895_30_fu_19950_p2;
wire   [0:0] or_ln895_15_fu_19956_p2;
wire   [0:0] xor_ln895_31_fu_19961_p2;
wire   [0:0] deleted_ones_15_fu_19940_p2;
wire   [0:0] xor_ln896_31_fu_19972_p2;
wire   [0:0] and_ln891_15_fu_19945_p2;
wire   [0:0] or_ln896_15_fu_19978_p2;
wire   [0:0] xor_ln896_258_fu_19984_p2;
wire   [0:0] overflow_15_fu_19966_p2;
wire   [0:0] underflow_15_fu_19990_p2;
wire   [0:0] or_ln346_15_fu_20003_p2;
wire   [31:0] select_ln346_30_fu_19995_p3;
wire  signed [31:0] sext_ln856_14_fu_19892_p1;
wire   [19:0] zext_ln377_16_fu_20020_p1;
wire  signed [19:0] sext_ln823_15_fu_20017_p1;
wire  signed [19:0] p_Val2_47_fu_20023_p2;
wire   [0:0] p_Result_48_fu_20033_p3;
wire   [0:0] xor_ln896_32_fu_20041_p2;
wire   [0:0] xor_ln888_29_fu_20052_p2;
wire   [0:0] or_ln888_16_fu_20057_p2;
wire   [0:0] tmp_93_fu_20068_p3;
wire   [0:0] xor_ln890_14_fu_20076_p2;
wire   [0:0] or_ln890_16_fu_20082_p2;
wire   [0:0] carry_30_fu_20047_p2;
wire   [0:0] deleted_zeros_13_fu_20063_p2;
wire   [0:0] xor_ln895_32_fu_20098_p2;
wire   [0:0] or_ln895_16_fu_20104_p2;
wire   [0:0] xor_ln895_33_fu_20110_p2;
wire   [0:0] deleted_ones_16_fu_20088_p2;
wire   [0:0] xor_ln896_33_fu_20121_p2;
wire   [0:0] and_ln891_16_fu_20093_p2;
wire   [0:0] or_ln896_16_fu_20127_p2;
wire   [0:0] xor_ln896_259_fu_20133_p2;
wire   [0:0] overflow_16_fu_20115_p2;
wire   [0:0] underflow_16_fu_20139_p2;
wire   [0:0] or_ln346_16_fu_20152_p2;
wire   [31:0] select_ln346_32_fu_20144_p3;
wire  signed [31:0] sext_ln856_15_fu_20029_p1;
wire   [21:0] zext_ln377_17_fu_20169_p1;
wire  signed [21:0] sext_ln823_16_fu_20166_p1;
wire  signed [21:0] p_Val2_50_fu_20172_p2;
wire   [0:0] p_Result_51_fu_20182_p3;
wire   [0:0] xor_ln896_34_fu_20190_p2;
wire   [0:0] xor_ln888_31_fu_20201_p2;
wire   [0:0] or_ln888_17_fu_20206_p2;
wire   [0:0] tmp_99_fu_20217_p3;
wire   [0:0] xor_ln890_15_fu_20225_p2;
wire   [0:0] or_ln890_17_fu_20231_p2;
wire   [0:0] carry_32_fu_20196_p2;
wire   [0:0] deleted_zeros_14_fu_20212_p2;
wire   [0:0] xor_ln895_34_fu_20247_p2;
wire   [0:0] or_ln895_17_fu_20253_p2;
wire   [0:0] xor_ln895_35_fu_20259_p2;
wire   [0:0] deleted_ones_17_fu_20237_p2;
wire   [0:0] xor_ln896_35_fu_20270_p2;
wire   [0:0] and_ln891_17_fu_20242_p2;
wire   [0:0] or_ln896_17_fu_20276_p2;
wire   [0:0] xor_ln896_260_fu_20282_p2;
wire   [0:0] overflow_17_fu_20264_p2;
wire   [0:0] underflow_17_fu_20288_p2;
wire   [0:0] or_ln346_17_fu_20301_p2;
wire   [31:0] select_ln346_34_fu_20293_p3;
wire  signed [31:0] sext_ln856_16_fu_20178_p1;
wire   [19:0] zext_ln377_18_fu_20318_p1;
wire  signed [19:0] sext_ln823_17_fu_20315_p1;
wire   [0:0] p_Result_54_fu_20327_p3;
wire   [0:0] xor_ln896_36_fu_20335_p2;
wire   [0:0] xor_ln888_33_fu_20346_p2;
wire   [0:0] or_ln888_18_fu_20351_p2;
wire   [0:0] tmp_105_fu_20362_p3;
wire   [0:0] xor_ln890_16_fu_20370_p2;
wire   [0:0] or_ln890_18_fu_20376_p2;
wire   [0:0] carry_34_fu_20341_p2;
wire   [0:0] deleted_zeros_15_fu_20357_p2;
wire   [0:0] xor_ln895_36_fu_20392_p2;
wire   [0:0] or_ln895_18_fu_20398_p2;
wire   [0:0] xor_ln895_37_fu_20404_p2;
wire   [0:0] deleted_ones_18_fu_20382_p2;
wire   [0:0] xor_ln896_37_fu_20415_p2;
wire   [0:0] and_ln891_18_fu_20387_p2;
wire   [0:0] or_ln896_18_fu_20421_p2;
wire   [0:0] xor_ln896_261_fu_20427_p2;
wire   [0:0] underflow_18_fu_20433_p2;
wire   [20:0] zext_ln377_19_fu_20447_p1;
wire  signed [20:0] sext_ln823_18_fu_20444_p1;
wire   [0:0] p_Result_57_fu_20456_p3;
wire   [0:0] xor_ln896_38_fu_20464_p2;
wire   [0:0] xor_ln888_35_fu_20475_p2;
wire   [0:0] or_ln888_19_fu_20480_p2;
wire   [0:0] tmp_111_fu_20491_p3;
wire   [0:0] xor_ln890_17_fu_20499_p2;
wire   [0:0] or_ln890_19_fu_20505_p2;
wire   [0:0] carry_36_fu_20470_p2;
wire   [0:0] deleted_zeros_16_fu_20486_p2;
wire   [0:0] xor_ln895_38_fu_20521_p2;
wire   [0:0] or_ln895_19_fu_20527_p2;
wire   [0:0] xor_ln895_39_fu_20533_p2;
wire   [0:0] deleted_ones_19_fu_20511_p2;
wire   [0:0] xor_ln896_39_fu_20544_p2;
wire   [0:0] and_ln891_19_fu_20516_p2;
wire   [0:0] or_ln896_19_fu_20550_p2;
wire   [0:0] xor_ln896_262_fu_20556_p2;
wire   [0:0] underflow_19_fu_20562_p2;
wire   [18:0] zext_ln377_20_fu_20576_p1;
wire  signed [18:0] sext_ln823_19_fu_20573_p1;
wire  signed [18:0] p_Val2_59_fu_20579_p2;
wire   [0:0] p_Result_60_fu_20589_p3;
wire   [0:0] xor_ln896_40_fu_20597_p2;
wire   [0:0] xor_ln888_37_fu_20608_p2;
wire   [0:0] or_ln888_20_fu_20613_p2;
wire   [0:0] tmp_117_fu_20624_p3;
wire   [0:0] xor_ln890_18_fu_20632_p2;
wire   [0:0] or_ln890_20_fu_20638_p2;
wire   [0:0] carry_38_fu_20603_p2;
wire   [0:0] deleted_zeros_17_fu_20619_p2;
wire   [0:0] xor_ln895_40_fu_20654_p2;
wire   [0:0] or_ln895_20_fu_20660_p2;
wire   [0:0] xor_ln895_41_fu_20666_p2;
wire   [0:0] deleted_ones_20_fu_20644_p2;
wire   [0:0] xor_ln896_41_fu_20677_p2;
wire   [0:0] and_ln891_20_fu_20649_p2;
wire   [0:0] or_ln896_20_fu_20683_p2;
wire   [0:0] xor_ln896_263_fu_20689_p2;
wire   [0:0] overflow_20_fu_20671_p2;
wire   [0:0] underflow_20_fu_20695_p2;
wire   [0:0] or_ln346_20_fu_20708_p2;
wire   [31:0] select_ln346_40_fu_20700_p3;
wire  signed [31:0] sext_ln856_19_fu_20585_p1;
wire   [19:0] zext_ln377_21_fu_20725_p1;
wire  signed [19:0] sext_ln823_20_fu_20722_p1;
wire   [0:0] p_Result_63_fu_20734_p3;
wire   [0:0] xor_ln896_42_fu_20742_p2;
wire   [0:0] xor_ln888_39_fu_20753_p2;
wire   [0:0] or_ln888_21_fu_20758_p2;
wire   [0:0] tmp_123_fu_20769_p3;
wire   [0:0] xor_ln890_19_fu_20777_p2;
wire   [0:0] or_ln890_21_fu_20783_p2;
wire   [0:0] carry_40_fu_20748_p2;
wire   [0:0] deleted_zeros_18_fu_20764_p2;
wire   [0:0] xor_ln895_42_fu_20799_p2;
wire   [0:0] or_ln895_21_fu_20805_p2;
wire   [0:0] xor_ln895_43_fu_20811_p2;
wire   [0:0] deleted_ones_21_fu_20789_p2;
wire   [0:0] xor_ln896_43_fu_20822_p2;
wire   [0:0] and_ln891_21_fu_20794_p2;
wire   [0:0] or_ln896_21_fu_20828_p2;
wire   [0:0] xor_ln896_264_fu_20834_p2;
wire   [0:0] underflow_21_fu_20840_p2;
wire   [19:0] zext_ln377_22_fu_20854_p1;
wire  signed [19:0] sext_ln823_21_fu_20851_p1;
wire   [0:0] p_Result_66_fu_20863_p3;
wire   [0:0] xor_ln896_44_fu_20871_p2;
wire   [0:0] xor_ln888_41_fu_20882_p2;
wire   [0:0] or_ln888_22_fu_20887_p2;
wire   [0:0] tmp_129_fu_20898_p3;
wire   [0:0] xor_ln890_20_fu_20906_p2;
wire   [0:0] or_ln890_22_fu_20912_p2;
wire   [0:0] carry_42_fu_20877_p2;
wire   [0:0] deleted_zeros_19_fu_20893_p2;
wire   [0:0] xor_ln895_44_fu_20928_p2;
wire   [0:0] or_ln895_22_fu_20934_p2;
wire   [0:0] xor_ln895_45_fu_20940_p2;
wire   [0:0] deleted_ones_22_fu_20918_p2;
wire   [0:0] xor_ln896_45_fu_20951_p2;
wire   [0:0] and_ln891_22_fu_20923_p2;
wire   [0:0] or_ln896_22_fu_20957_p2;
wire   [0:0] xor_ln896_265_fu_20963_p2;
wire   [0:0] underflow_22_fu_20969_p2;
wire   [14:0] zext_ln377_23_fu_20983_p1;
wire  signed [14:0] sext_ln823_22_fu_20980_p1;
wire   [0:0] p_Result_69_fu_20992_p3;
wire   [0:0] xor_ln896_46_fu_21000_p2;
wire   [0:0] xor_ln888_43_fu_21011_p2;
wire   [0:0] or_ln888_23_fu_21016_p2;
wire   [0:0] tmp_135_fu_21027_p3;
wire   [0:0] xor_ln890_21_fu_21035_p2;
wire   [0:0] or_ln890_23_fu_21041_p2;
wire   [0:0] carry_44_fu_21006_p2;
wire   [0:0] deleted_zeros_20_fu_21022_p2;
wire   [0:0] xor_ln895_46_fu_21057_p2;
wire   [0:0] or_ln895_23_fu_21063_p2;
wire   [0:0] xor_ln895_47_fu_21069_p2;
wire   [0:0] deleted_ones_23_fu_21047_p2;
wire   [0:0] xor_ln896_47_fu_21080_p2;
wire   [0:0] and_ln891_23_fu_21052_p2;
wire   [0:0] or_ln896_23_fu_21086_p2;
wire   [0:0] xor_ln896_266_fu_21092_p2;
wire   [0:0] underflow_23_fu_21098_p2;
wire   [31:0] select_ln346_48_fu_21112_p3;
wire  signed [31:0] sext_ln856_23_fu_21109_p1;
wire   [21:0] zext_ln377_25_fu_21129_p1;
wire  signed [21:0] sext_ln823_24_fu_21126_p1;
wire   [0:0] p_Result_75_fu_21138_p3;
wire   [0:0] xor_ln896_50_fu_21146_p2;
wire   [0:0] xor_ln888_47_fu_21157_p2;
wire   [0:0] or_ln888_25_fu_21162_p2;
wire   [0:0] tmp_147_fu_21173_p3;
wire   [0:0] xor_ln890_23_fu_21181_p2;
wire   [0:0] or_ln890_25_fu_21187_p2;
wire   [0:0] carry_48_fu_21152_p2;
wire   [0:0] deleted_zeros_22_fu_21168_p2;
wire   [0:0] xor_ln895_50_fu_21203_p2;
wire   [0:0] or_ln895_25_fu_21209_p2;
wire   [0:0] xor_ln895_51_fu_21215_p2;
wire   [0:0] deleted_ones_25_fu_21193_p2;
wire   [0:0] xor_ln896_51_fu_21226_p2;
wire   [0:0] and_ln891_25_fu_21198_p2;
wire   [0:0] or_ln896_25_fu_21232_p2;
wire   [0:0] xor_ln896_268_fu_21238_p2;
wire   [0:0] underflow_25_fu_21244_p2;
wire   [19:0] zext_ln377_26_fu_21258_p1;
wire  signed [19:0] sext_ln823_25_fu_21255_p1;
wire   [0:0] p_Result_78_fu_21267_p3;
wire   [0:0] xor_ln896_52_fu_21275_p2;
wire   [0:0] xor_ln888_49_fu_21286_p2;
wire   [0:0] or_ln888_26_fu_21291_p2;
wire   [0:0] tmp_153_fu_21302_p3;
wire   [0:0] xor_ln890_24_fu_21310_p2;
wire   [0:0] or_ln890_26_fu_21316_p2;
wire   [0:0] carry_50_fu_21281_p2;
wire   [0:0] deleted_zeros_23_fu_21297_p2;
wire   [0:0] xor_ln895_52_fu_21332_p2;
wire   [0:0] or_ln895_26_fu_21338_p2;
wire   [0:0] xor_ln895_53_fu_21344_p2;
wire   [0:0] deleted_ones_26_fu_21322_p2;
wire   [0:0] xor_ln896_53_fu_21355_p2;
wire   [0:0] and_ln891_26_fu_21327_p2;
wire   [0:0] or_ln896_26_fu_21361_p2;
wire   [0:0] xor_ln896_269_fu_21367_p2;
wire   [0:0] underflow_26_fu_21373_p2;
wire   [0:0] tmp_156_fu_21434_p3;
wire   [31:0] zext_ln377_27_fu_21442_p1;
wire   [31:0] p_Val2_79_fu_21416_p4;
wire   [19:0] p_Val2_82_fu_21476_p4;
wire   [0:0] tmp_162_fu_21498_p3;
wire   [20:0] zext_ln377_28_fu_21506_p1;
wire  signed [20:0] sext_ln823_26_fu_21486_p1;
wire   [18:0] p_Val2_85_fu_21540_p4;
wire   [0:0] tmp_168_fu_21562_p3;
wire   [19:0] zext_ln377_29_fu_21570_p1;
wire  signed [19:0] sext_ln823_27_fu_21550_p1;
wire   [19:0] p_Val2_88_fu_21604_p4;
wire   [0:0] tmp_174_fu_21626_p3;
wire   [20:0] zext_ln377_30_fu_21634_p1;
wire  signed [20:0] sext_ln823_28_fu_21614_p1;
wire   [18:0] p_Val2_91_fu_21668_p4;
wire   [0:0] tmp_180_fu_21690_p3;
wire   [19:0] zext_ln377_31_fu_21698_p1;
wire  signed [19:0] sext_ln823_29_fu_21678_p1;
wire   [16:0] p_Val2_94_fu_21732_p4;
wire   [0:0] tmp_186_fu_21754_p3;
wire   [17:0] zext_ln377_32_fu_21762_p1;
wire  signed [17:0] sext_ln823_30_fu_21742_p1;
wire   [16:0] p_Val2_97_fu_21796_p4;
wire   [0:0] tmp_192_fu_21818_p3;
wire   [17:0] zext_ln377_33_fu_21826_p1;
wire  signed [17:0] sext_ln823_31_fu_21806_p1;
wire   [21:0] p_Val2_100_fu_21860_p4;
wire   [0:0] tmp_198_fu_21882_p3;
wire   [22:0] zext_ln377_34_fu_21890_p1;
wire  signed [22:0] sext_ln823_32_fu_21870_p1;
wire   [0:0] tmp_204_fu_21942_p3;
wire   [31:0] zext_ln377_35_fu_21950_p1;
wire   [31:0] p_Val2_103_fu_21924_p4;
wire   [36:0] shl_ln1273_3_fu_22131_p3;
wire  signed [37:0] sext_ln1273_3_fu_22138_p1;
wire  signed [37:0] sext_ln70_22_fu_21989_p1;
wire   [37:0] r_V_36_fu_22142_p2;
wire   [13:0] p_Val2_115_fu_22156_p4;
wire   [0:0] tmp_228_fu_22178_p3;
wire   [14:0] zext_ln377_39_fu_22186_p1;
wire  signed [14:0] sext_ln823_36_fu_22166_p1;
wire   [0:0] p_Result_117_fu_22196_p3;
wire   [0:0] p_Result_116_fu_22170_p3;
wire   [0:0] xor_ln896_78_fu_22204_p2;
wire   [0:0] xor_ln888_75_fu_22224_p2;
wire   [0:0] Range2_all_ones_37_fu_22216_p3;
wire   [0:0] or_ln888_39_fu_22230_p2;
wire   [0:0] tmp_231_fu_22242_p3;
wire   [0:0] xor_ln890_37_fu_22250_p2;
wire   [0:0] or_ln890_39_fu_22256_p2;
wire   [0:0] carry_76_fu_22210_p2;
wire   [0:0] deleted_zeros_36_fu_22236_p2;
wire   [0:0] xor_ln895_78_fu_22274_p2;
wire   [0:0] p_Result_115_fu_22148_p3;
wire   [0:0] or_ln895_39_fu_22280_p2;
wire   [0:0] xor_ln895_79_fu_22286_p2;
wire   [0:0] deleted_ones_39_fu_22262_p2;
wire   [0:0] xor_ln896_79_fu_22298_p2;
wire   [0:0] and_ln891_39_fu_22268_p2;
wire   [0:0] or_ln896_39_fu_22304_p2;
wire   [0:0] xor_ln896_282_fu_22310_p2;
wire   [0:0] underflow_39_fu_22316_p2;
wire  signed [31:0] rhs_fu_18606_p3;
wire  signed [32:0] sext_ln813_fu_22538_p1;
wire   [32:0] ret_V_fu_22542_p2;
wire   [31:0] p_Val2_241_fu_22556_p2;
wire   [0:0] p_Result_241_fu_22548_p3;
wire   [0:0] p_Result_242_fu_22562_p3;
wire   [0:0] xor_ln895_162_fu_22570_p2;
wire   [0:0] xor_ln896_162_fu_22582_p2;
wire   [0:0] xor_ln302_fu_22594_p2;
wire   [0:0] overflow_81_fu_22576_p2;
wire   [0:0] xor_ln302_1_fu_22600_p2;
wire   [0:0] underflow_81_fu_22588_p2;
wire   [0:0] or_ln302_fu_22606_p2;
wire   [31:0] select_ln302_fu_22612_p3;
wire   [31:0] select_ln350_fu_22620_p3;
wire  signed [31:0] rhs_1_fu_18731_p3;
wire  signed [32:0] sext_ln813_1_fu_22636_p1;
wire   [32:0] ret_V_1_fu_22640_p2;
wire   [31:0] p_Val2_243_fu_22654_p2;
wire   [0:0] p_Result_243_fu_22646_p3;
wire   [0:0] p_Result_244_fu_22660_p3;
wire   [0:0] xor_ln895_163_fu_22668_p2;
wire   [0:0] xor_ln896_163_fu_22680_p2;
wire   [0:0] xor_ln302_2_fu_22692_p2;
wire   [0:0] overflow_82_fu_22674_p2;
wire   [0:0] xor_ln302_3_fu_22698_p2;
wire   [0:0] underflow_82_fu_22686_p2;
wire   [0:0] or_ln302_1_fu_22704_p2;
wire   [31:0] select_ln302_2_fu_22710_p3;
wire   [31:0] select_ln350_1_fu_22718_p3;
wire  signed [31:0] rhs_2_fu_18749_p3;
wire  signed [32:0] sext_ln813_2_fu_22734_p1;
wire   [32:0] ret_V_2_fu_22738_p2;
wire   [31:0] p_Val2_245_fu_22752_p2;
wire   [0:0] p_Result_245_fu_22744_p3;
wire   [0:0] p_Result_246_fu_22758_p3;
wire   [0:0] xor_ln895_164_fu_22766_p2;
wire   [0:0] xor_ln896_164_fu_22778_p2;
wire   [0:0] xor_ln302_4_fu_22790_p2;
wire   [0:0] overflow_83_fu_22772_p2;
wire   [0:0] xor_ln302_5_fu_22796_p2;
wire   [0:0] underflow_83_fu_22784_p2;
wire   [0:0] or_ln302_2_fu_22802_p2;
wire   [31:0] select_ln302_4_fu_22808_p3;
wire   [31:0] select_ln350_2_fu_22816_p3;
wire  signed [31:0] rhs_3_fu_18873_p3;
wire  signed [32:0] sext_ln813_3_fu_22832_p1;
wire   [32:0] ret_V_3_fu_22836_p2;
wire   [31:0] p_Val2_247_fu_22850_p2;
wire   [0:0] p_Result_247_fu_22842_p3;
wire   [0:0] p_Result_248_fu_22856_p3;
wire   [0:0] xor_ln895_165_fu_22864_p2;
wire   [0:0] xor_ln896_165_fu_22876_p2;
wire   [0:0] xor_ln302_6_fu_22888_p2;
wire   [0:0] overflow_84_fu_22870_p2;
wire   [0:0] xor_ln302_7_fu_22894_p2;
wire   [0:0] underflow_84_fu_22882_p2;
wire   [0:0] or_ln302_3_fu_22900_p2;
wire   [31:0] select_ln302_6_fu_22906_p3;
wire   [31:0] select_ln350_3_fu_22914_p3;
wire  signed [31:0] rhs_4_fu_18998_p3;
wire  signed [32:0] sext_ln813_4_fu_22930_p1;
wire   [32:0] ret_V_4_fu_22934_p2;
wire   [31:0] p_Val2_249_fu_22948_p2;
wire   [0:0] p_Result_249_fu_22940_p3;
wire   [0:0] p_Result_250_fu_22954_p3;
wire   [0:0] xor_ln895_166_fu_22962_p2;
wire   [0:0] xor_ln896_166_fu_22974_p2;
wire   [0:0] xor_ln302_8_fu_22986_p2;
wire   [0:0] overflow_85_fu_22968_p2;
wire   [0:0] xor_ln302_9_fu_22992_p2;
wire   [0:0] underflow_85_fu_22980_p2;
wire   [0:0] or_ln302_4_fu_22998_p2;
wire   [31:0] select_ln302_8_fu_23004_p3;
wire   [31:0] select_ln350_4_fu_23012_p3;
wire  signed [31:0] rhs_5_fu_19123_p3;
wire  signed [32:0] sext_ln813_5_fu_23028_p1;
wire   [32:0] ret_V_5_fu_23032_p2;
wire   [31:0] p_Val2_251_fu_23046_p2;
wire   [0:0] p_Result_251_fu_23038_p3;
wire   [0:0] p_Result_252_fu_23052_p3;
wire   [0:0] xor_ln895_167_fu_23060_p2;
wire   [0:0] xor_ln896_167_fu_23072_p2;
wire   [0:0] xor_ln302_10_fu_23084_p2;
wire   [0:0] overflow_86_fu_23066_p2;
wire   [0:0] xor_ln302_11_fu_23090_p2;
wire   [0:0] underflow_86_fu_23078_p2;
wire   [0:0] or_ln302_5_fu_23096_p2;
wire   [31:0] select_ln302_10_fu_23102_p3;
wire   [31:0] select_ln350_5_fu_23110_p3;
wire  signed [31:0] rhs_6_fu_19141_p3;
wire  signed [32:0] sext_ln813_6_fu_23126_p1;
wire   [32:0] ret_V_6_fu_23130_p2;
wire   [31:0] p_Val2_253_fu_23144_p2;
wire   [0:0] p_Result_253_fu_23136_p3;
wire   [0:0] p_Result_254_fu_23150_p3;
wire   [0:0] xor_ln895_168_fu_23158_p2;
wire   [0:0] xor_ln896_168_fu_23170_p2;
wire   [0:0] xor_ln302_12_fu_23182_p2;
wire   [0:0] overflow_87_fu_23164_p2;
wire   [0:0] xor_ln302_13_fu_23188_p2;
wire   [0:0] underflow_87_fu_23176_p2;
wire   [0:0] or_ln302_6_fu_23194_p2;
wire   [31:0] select_ln302_12_fu_23200_p3;
wire   [31:0] select_ln350_6_fu_23208_p3;
wire  signed [31:0] rhs_7_fu_19262_p3;
wire  signed [32:0] sext_ln813_7_fu_23224_p1;
wire   [32:0] ret_V_7_fu_23228_p2;
wire   [31:0] p_Val2_255_fu_23242_p2;
wire   [0:0] p_Result_255_fu_23234_p3;
wire   [0:0] p_Result_256_fu_23248_p3;
wire   [0:0] xor_ln895_169_fu_23256_p2;
wire   [0:0] xor_ln896_169_fu_23268_p2;
wire   [0:0] xor_ln302_14_fu_23280_p2;
wire   [0:0] overflow_88_fu_23262_p2;
wire   [0:0] xor_ln302_15_fu_23286_p2;
wire   [0:0] underflow_88_fu_23274_p2;
wire   [0:0] or_ln302_7_fu_23292_p2;
wire   [31:0] select_ln302_14_fu_23298_p3;
wire   [31:0] select_ln350_7_fu_23306_p3;
wire  signed [31:0] rhs_8_fu_19386_p3;
wire  signed [32:0] sext_ln813_8_fu_23322_p1;
wire   [32:0] ret_V_8_fu_23326_p2;
wire   [31:0] p_Val2_257_fu_23340_p2;
wire   [0:0] p_Result_257_fu_23332_p3;
wire   [0:0] p_Result_258_fu_23346_p3;
wire   [0:0] xor_ln895_170_fu_23354_p2;
wire   [0:0] xor_ln896_170_fu_23366_p2;
wire   [0:0] xor_ln302_16_fu_23378_p2;
wire   [0:0] overflow_89_fu_23360_p2;
wire   [0:0] xor_ln302_17_fu_23384_p2;
wire   [0:0] underflow_89_fu_23372_p2;
wire   [0:0] or_ln302_8_fu_23390_p2;
wire   [31:0] select_ln302_16_fu_23396_p3;
wire   [31:0] select_ln350_8_fu_23404_p3;
wire  signed [31:0] lhs_fu_22628_p3;
wire  signed [31:0] rhs_9_fu_19535_p3;
wire  signed [32:0] sext_ln813_10_fu_23424_p1;
wire  signed [32:0] sext_ln813_9_fu_23420_p1;
wire   [32:0] ret_V_9_fu_23428_p2;
wire   [31:0] p_Val2_259_fu_23442_p2;
wire   [0:0] p_Result_259_fu_23434_p3;
wire   [0:0] p_Result_260_fu_23448_p3;
wire   [0:0] xor_ln895_171_fu_23456_p2;
wire   [0:0] xor_ln896_171_fu_23468_p2;
wire   [0:0] xor_ln302_18_fu_23480_p2;
wire   [0:0] overflow_90_fu_23462_p2;
wire   [0:0] xor_ln302_19_fu_23486_p2;
wire   [0:0] underflow_90_fu_23474_p2;
wire   [0:0] or_ln302_9_fu_23492_p2;
wire   [31:0] select_ln302_18_fu_23498_p3;
wire   [31:0] select_ln350_9_fu_23506_p3;
wire  signed [31:0] lhs_1_fu_22726_p3;
wire  signed [31:0] rhs_10_fu_19553_p3;
wire  signed [32:0] sext_ln813_12_fu_23526_p1;
wire  signed [32:0] sext_ln813_11_fu_23522_p1;
wire   [32:0] ret_V_10_fu_23530_p2;
wire   [31:0] p_Val2_261_fu_23544_p2;
wire   [0:0] p_Result_261_fu_23536_p3;
wire   [0:0] p_Result_262_fu_23550_p3;
wire   [0:0] xor_ln895_172_fu_23558_p2;
wire   [0:0] xor_ln896_172_fu_23570_p2;
wire   [0:0] xor_ln302_20_fu_23582_p2;
wire   [0:0] overflow_91_fu_23564_p2;
wire   [0:0] xor_ln302_21_fu_23588_p2;
wire   [0:0] underflow_91_fu_23576_p2;
wire   [0:0] or_ln302_10_fu_23594_p2;
wire   [31:0] select_ln302_20_fu_23600_p3;
wire   [31:0] select_ln350_10_fu_23608_p3;
wire  signed [31:0] lhs_2_fu_22824_p3;
wire  signed [31:0] rhs_11_fu_19570_p3;
wire  signed [32:0] sext_ln813_14_fu_23628_p1;
wire  signed [32:0] sext_ln813_13_fu_23624_p1;
wire   [32:0] ret_V_11_fu_23632_p2;
wire   [31:0] p_Val2_263_fu_23646_p2;
wire   [0:0] p_Result_263_fu_23638_p3;
wire   [0:0] p_Result_264_fu_23652_p3;
wire   [0:0] xor_ln895_173_fu_23660_p2;
wire   [0:0] xor_ln896_173_fu_23672_p2;
wire   [0:0] xor_ln302_22_fu_23684_p2;
wire   [0:0] overflow_92_fu_23666_p2;
wire   [0:0] xor_ln302_23_fu_23690_p2;
wire   [0:0] underflow_92_fu_23678_p2;
wire   [0:0] or_ln302_11_fu_23696_p2;
wire   [31:0] select_ln302_22_fu_23702_p3;
wire   [31:0] select_ln350_11_fu_23710_p3;
wire  signed [31:0] lhs_3_fu_22922_p3;
wire  signed [31:0] rhs_12_fu_19718_p3;
wire  signed [32:0] sext_ln813_16_fu_23730_p1;
wire  signed [32:0] sext_ln813_15_fu_23726_p1;
wire   [32:0] ret_V_12_fu_23734_p2;
wire   [31:0] p_Val2_265_fu_23748_p2;
wire   [0:0] p_Result_265_fu_23740_p3;
wire   [0:0] p_Result_266_fu_23754_p3;
wire   [0:0] xor_ln895_174_fu_23762_p2;
wire   [0:0] xor_ln896_174_fu_23774_p2;
wire   [0:0] xor_ln302_24_fu_23786_p2;
wire   [0:0] overflow_93_fu_23768_p2;
wire   [0:0] xor_ln302_25_fu_23792_p2;
wire   [0:0] underflow_93_fu_23780_p2;
wire   [0:0] or_ln302_12_fu_23798_p2;
wire   [31:0] select_ln302_24_fu_23804_p3;
wire   [31:0] select_ln350_12_fu_23812_p3;
wire  signed [31:0] lhs_4_fu_23020_p3;
wire  signed [31:0] rhs_13_fu_19867_p3;
wire  signed [32:0] sext_ln813_18_fu_23832_p1;
wire  signed [32:0] sext_ln813_17_fu_23828_p1;
wire   [32:0] ret_V_13_fu_23836_p2;
wire   [31:0] p_Val2_267_fu_23850_p2;
wire   [0:0] p_Result_267_fu_23842_p3;
wire   [0:0] p_Result_268_fu_23856_p3;
wire   [0:0] xor_ln895_175_fu_23864_p2;
wire   [0:0] xor_ln896_175_fu_23876_p2;
wire   [0:0] xor_ln302_26_fu_23888_p2;
wire   [0:0] overflow_94_fu_23870_p2;
wire   [0:0] xor_ln302_27_fu_23894_p2;
wire   [0:0] underflow_94_fu_23882_p2;
wire   [0:0] or_ln302_13_fu_23900_p2;
wire   [31:0] select_ln302_26_fu_23906_p3;
wire   [31:0] select_ln350_13_fu_23914_p3;
wire  signed [31:0] lhs_5_fu_23118_p3;
wire  signed [31:0] rhs_14_fu_19885_p3;
wire  signed [32:0] sext_ln813_20_fu_23934_p1;
wire  signed [32:0] sext_ln813_19_fu_23930_p1;
wire   [32:0] ret_V_14_fu_23938_p2;
wire   [31:0] p_Val2_269_fu_23952_p2;
wire   [0:0] p_Result_269_fu_23944_p3;
wire   [0:0] p_Result_270_fu_23958_p3;
wire   [0:0] xor_ln895_176_fu_23966_p2;
wire   [0:0] xor_ln896_176_fu_23978_p2;
wire   [0:0] xor_ln302_28_fu_23990_p2;
wire   [0:0] overflow_95_fu_23972_p2;
wire   [0:0] xor_ln302_29_fu_23996_p2;
wire   [0:0] underflow_95_fu_23984_p2;
wire   [0:0] or_ln302_14_fu_24002_p2;
wire   [31:0] select_ln302_28_fu_24008_p3;
wire   [31:0] select_ln350_14_fu_24016_p3;
wire  signed [31:0] lhs_6_fu_23216_p3;
wire  signed [31:0] rhs_15_fu_20009_p3;
wire  signed [32:0] sext_ln813_22_fu_24036_p1;
wire  signed [32:0] sext_ln813_21_fu_24032_p1;
wire   [32:0] ret_V_15_fu_24040_p2;
wire   [31:0] p_Val2_271_fu_24054_p2;
wire   [0:0] p_Result_271_fu_24046_p3;
wire   [0:0] p_Result_272_fu_24060_p3;
wire   [0:0] xor_ln895_177_fu_24068_p2;
wire   [0:0] xor_ln896_177_fu_24080_p2;
wire   [0:0] xor_ln302_30_fu_24092_p2;
wire   [0:0] overflow_96_fu_24074_p2;
wire   [0:0] xor_ln302_31_fu_24098_p2;
wire   [0:0] underflow_96_fu_24086_p2;
wire   [0:0] or_ln302_15_fu_24104_p2;
wire   [31:0] select_ln302_30_fu_24110_p3;
wire   [31:0] select_ln350_15_fu_24118_p3;
wire  signed [31:0] lhs_7_fu_23314_p3;
wire  signed [31:0] rhs_16_fu_20158_p3;
wire  signed [32:0] sext_ln813_24_fu_24138_p1;
wire  signed [32:0] sext_ln813_23_fu_24134_p1;
wire   [32:0] ret_V_16_fu_24142_p2;
wire   [31:0] p_Val2_273_fu_24156_p2;
wire   [0:0] p_Result_273_fu_24148_p3;
wire   [0:0] p_Result_274_fu_24162_p3;
wire   [0:0] xor_ln895_178_fu_24170_p2;
wire   [0:0] xor_ln896_178_fu_24182_p2;
wire   [0:0] xor_ln302_32_fu_24194_p2;
wire   [0:0] overflow_97_fu_24176_p2;
wire   [0:0] xor_ln302_33_fu_24200_p2;
wire   [0:0] underflow_97_fu_24188_p2;
wire   [0:0] or_ln302_16_fu_24206_p2;
wire   [31:0] select_ln302_32_fu_24212_p3;
wire   [31:0] select_ln350_16_fu_24220_p3;
wire  signed [31:0] lhs_8_fu_23412_p3;
wire  signed [31:0] rhs_17_fu_20307_p3;
wire  signed [32:0] sext_ln813_26_fu_24240_p1;
wire  signed [32:0] sext_ln813_25_fu_24236_p1;
wire   [32:0] ret_V_17_fu_24244_p2;
wire   [31:0] p_Val2_275_fu_24258_p2;
wire   [0:0] p_Result_275_fu_24250_p3;
wire   [0:0] p_Result_276_fu_24264_p3;
wire   [0:0] xor_ln895_179_fu_24272_p2;
wire   [0:0] xor_ln896_179_fu_24284_p2;
wire   [0:0] xor_ln302_34_fu_24296_p2;
wire   [0:0] overflow_98_fu_24278_p2;
wire   [0:0] xor_ln302_35_fu_24302_p2;
wire   [0:0] underflow_98_fu_24290_p2;
wire   [0:0] or_ln302_17_fu_24308_p2;
wire   [31:0] select_ln302_34_fu_24314_p3;
wire   [31:0] select_ln350_17_fu_24322_p3;
wire  signed [31:0] lhs_11_fu_23718_p3;
wire  signed [31:0] rhs_20_fu_20714_p3;
wire  signed [32:0] sext_ln813_32_fu_24342_p1;
wire  signed [32:0] sext_ln813_31_fu_24338_p1;
wire   [32:0] ret_V_20_fu_24346_p2;
wire  signed [31:0] lhs_15_fu_24126_p3;
wire  signed [31:0] rhs_24_fu_21119_p3;
wire  signed [32:0] sext_ln813_40_fu_24378_p1;
wire  signed [32:0] sext_ln813_39_fu_24374_p1;
wire   [32:0] ret_V_24_fu_24382_p2;
wire   [31:0] select_ln346_36_fu_24413_p3;
wire  signed [31:0] sext_ln856_17_fu_24410_p1;
wire   [31:0] select_ln346_38_fu_24430_p3;
wire  signed [31:0] sext_ln856_18_fu_24427_p1;
wire   [31:0] select_ln346_42_fu_24447_p3;
wire  signed [31:0] sext_ln856_20_fu_24444_p1;
wire   [31:0] select_ln346_44_fu_24464_p3;
wire  signed [31:0] sext_ln856_21_fu_24461_p1;
wire   [31:0] select_ln346_46_fu_24481_p3;
wire  signed [31:0] sext_ln856_22_fu_24478_p1;
wire   [31:0] select_ln346_50_fu_24498_p3;
wire  signed [31:0] sext_ln856_24_fu_24495_p1;
wire   [31:0] select_ln346_52_fu_24515_p3;
wire  signed [31:0] sext_ln856_25_fu_24512_p1;
wire   [0:0] xor_ln896_54_fu_24529_p2;
wire   [0:0] xor_ln888_51_fu_24539_p2;
wire   [0:0] or_ln888_27_fu_24544_p2;
wire   [0:0] tmp_159_fu_24554_p3;
wire   [0:0] xor_ln890_25_fu_24562_p2;
wire   [0:0] or_ln890_27_fu_24568_p2;
wire   [0:0] carry_52_fu_24534_p2;
wire   [0:0] deleted_zeros_24_fu_24549_p2;
wire   [0:0] xor_ln895_54_fu_24584_p2;
wire   [0:0] or_ln895_27_fu_24590_p2;
wire   [0:0] xor_ln895_55_fu_24595_p2;
wire   [0:0] deleted_ones_27_fu_24574_p2;
wire   [0:0] xor_ln896_55_fu_24606_p2;
wire   [0:0] and_ln891_27_fu_24579_p2;
wire   [0:0] or_ln896_27_fu_24612_p2;
wire   [0:0] xor_ln896_270_fu_24618_p2;
wire   [0:0] overflow_27_fu_24600_p2;
wire   [0:0] underflow_27_fu_24624_p2;
wire   [0:0] or_ln346_27_fu_24637_p2;
wire   [31:0] select_ln346_54_fu_24629_p3;
wire   [0:0] xor_ln896_56_fu_24653_p2;
wire   [0:0] xor_ln888_53_fu_24663_p2;
wire   [0:0] or_ln888_28_fu_24668_p2;
wire   [0:0] tmp_165_fu_24678_p3;
wire   [0:0] xor_ln890_26_fu_24686_p2;
wire   [0:0] or_ln890_28_fu_24692_p2;
wire   [0:0] carry_54_fu_24658_p2;
wire   [0:0] deleted_zeros_25_fu_24673_p2;
wire   [0:0] xor_ln895_56_fu_24708_p2;
wire   [0:0] or_ln895_28_fu_24714_p2;
wire   [0:0] xor_ln895_57_fu_24719_p2;
wire   [0:0] deleted_ones_28_fu_24698_p2;
wire   [0:0] xor_ln896_57_fu_24730_p2;
wire   [0:0] and_ln891_28_fu_24703_p2;
wire   [0:0] or_ln896_28_fu_24736_p2;
wire   [0:0] xor_ln896_271_fu_24742_p2;
wire   [0:0] overflow_28_fu_24724_p2;
wire   [0:0] underflow_28_fu_24748_p2;
wire   [0:0] or_ln346_28_fu_24761_p2;
wire   [31:0] select_ln346_56_fu_24753_p3;
wire  signed [31:0] sext_ln856_26_fu_24650_p1;
wire   [0:0] xor_ln896_58_fu_24778_p2;
wire   [0:0] xor_ln888_55_fu_24788_p2;
wire   [0:0] or_ln888_29_fu_24793_p2;
wire   [0:0] tmp_171_fu_24803_p3;
wire   [0:0] xor_ln890_27_fu_24811_p2;
wire   [0:0] or_ln890_29_fu_24817_p2;
wire   [0:0] carry_56_fu_24783_p2;
wire   [0:0] deleted_zeros_26_fu_24798_p2;
wire   [0:0] xor_ln895_58_fu_24833_p2;
wire   [0:0] or_ln895_29_fu_24839_p2;
wire   [0:0] xor_ln895_59_fu_24844_p2;
wire   [0:0] deleted_ones_29_fu_24823_p2;
wire   [0:0] xor_ln896_59_fu_24855_p2;
wire   [0:0] and_ln891_29_fu_24828_p2;
wire   [0:0] or_ln896_29_fu_24861_p2;
wire   [0:0] xor_ln896_272_fu_24867_p2;
wire   [0:0] overflow_29_fu_24849_p2;
wire   [0:0] underflow_29_fu_24873_p2;
wire   [0:0] or_ln346_29_fu_24886_p2;
wire   [31:0] select_ln346_58_fu_24878_p3;
wire  signed [31:0] sext_ln856_27_fu_24775_p1;
wire   [0:0] xor_ln896_60_fu_24903_p2;
wire   [0:0] xor_ln888_57_fu_24913_p2;
wire   [0:0] or_ln888_30_fu_24918_p2;
wire   [0:0] tmp_177_fu_24928_p3;
wire   [0:0] xor_ln890_28_fu_24936_p2;
wire   [0:0] or_ln890_30_fu_24942_p2;
wire   [0:0] carry_58_fu_24908_p2;
wire   [0:0] deleted_zeros_27_fu_24923_p2;
wire   [0:0] xor_ln895_60_fu_24958_p2;
wire   [0:0] or_ln895_30_fu_24964_p2;
wire   [0:0] xor_ln895_61_fu_24969_p2;
wire   [0:0] deleted_ones_30_fu_24948_p2;
wire   [0:0] xor_ln896_61_fu_24980_p2;
wire   [0:0] and_ln891_30_fu_24953_p2;
wire   [0:0] or_ln896_30_fu_24986_p2;
wire   [0:0] xor_ln896_273_fu_24992_p2;
wire   [0:0] overflow_30_fu_24974_p2;
wire   [0:0] underflow_30_fu_24998_p2;
wire   [0:0] or_ln346_30_fu_25011_p2;
wire   [31:0] select_ln346_60_fu_25003_p3;
wire  signed [31:0] sext_ln856_28_fu_24900_p1;
wire   [0:0] xor_ln896_62_fu_25028_p2;
wire   [0:0] xor_ln888_59_fu_25038_p2;
wire   [0:0] or_ln888_31_fu_25043_p2;
wire   [0:0] tmp_183_fu_25053_p3;
wire   [0:0] xor_ln890_29_fu_25061_p2;
wire   [0:0] or_ln890_31_fu_25067_p2;
wire   [0:0] carry_60_fu_25033_p2;
wire   [0:0] deleted_zeros_28_fu_25048_p2;
wire   [0:0] xor_ln895_62_fu_25083_p2;
wire   [0:0] or_ln895_31_fu_25089_p2;
wire   [0:0] xor_ln895_63_fu_25094_p2;
wire   [0:0] deleted_ones_31_fu_25073_p2;
wire   [0:0] xor_ln896_63_fu_25105_p2;
wire   [0:0] and_ln891_31_fu_25078_p2;
wire   [0:0] or_ln896_31_fu_25111_p2;
wire   [0:0] xor_ln896_274_fu_25117_p2;
wire   [0:0] overflow_31_fu_25099_p2;
wire   [0:0] underflow_31_fu_25123_p2;
wire   [0:0] or_ln346_31_fu_25136_p2;
wire   [31:0] select_ln346_62_fu_25128_p3;
wire  signed [31:0] sext_ln856_29_fu_25025_p1;
wire   [0:0] xor_ln896_64_fu_25153_p2;
wire   [0:0] xor_ln888_61_fu_25163_p2;
wire   [0:0] or_ln888_32_fu_25168_p2;
wire   [0:0] tmp_189_fu_25178_p3;
wire   [0:0] xor_ln890_30_fu_25186_p2;
wire   [0:0] or_ln890_32_fu_25192_p2;
wire   [0:0] carry_62_fu_25158_p2;
wire   [0:0] deleted_zeros_29_fu_25173_p2;
wire   [0:0] xor_ln895_64_fu_25208_p2;
wire   [0:0] or_ln895_32_fu_25214_p2;
wire   [0:0] xor_ln895_65_fu_25219_p2;
wire   [0:0] deleted_ones_32_fu_25198_p2;
wire   [0:0] xor_ln896_65_fu_25230_p2;
wire   [0:0] and_ln891_32_fu_25203_p2;
wire   [0:0] or_ln896_32_fu_25236_p2;
wire   [0:0] xor_ln896_275_fu_25242_p2;
wire   [0:0] overflow_32_fu_25224_p2;
wire   [0:0] underflow_32_fu_25248_p2;
wire   [0:0] or_ln346_32_fu_25261_p2;
wire   [31:0] select_ln346_64_fu_25253_p3;
wire  signed [31:0] sext_ln856_30_fu_25150_p1;
wire   [0:0] xor_ln896_66_fu_25278_p2;
wire   [0:0] xor_ln888_63_fu_25288_p2;
wire   [0:0] or_ln888_33_fu_25293_p2;
wire   [0:0] tmp_195_fu_25303_p3;
wire   [0:0] xor_ln890_31_fu_25311_p2;
wire   [0:0] or_ln890_33_fu_25317_p2;
wire   [0:0] carry_64_fu_25283_p2;
wire   [0:0] deleted_zeros_30_fu_25298_p2;
wire   [0:0] xor_ln895_66_fu_25333_p2;
wire   [0:0] or_ln895_33_fu_25339_p2;
wire   [0:0] xor_ln895_67_fu_25344_p2;
wire   [0:0] deleted_ones_33_fu_25323_p2;
wire   [0:0] xor_ln896_67_fu_25355_p2;
wire   [0:0] and_ln891_33_fu_25328_p2;
wire   [0:0] or_ln896_33_fu_25361_p2;
wire   [0:0] xor_ln896_276_fu_25367_p2;
wire   [0:0] overflow_33_fu_25349_p2;
wire   [0:0] underflow_33_fu_25373_p2;
wire   [0:0] or_ln346_33_fu_25386_p2;
wire   [31:0] select_ln346_66_fu_25378_p3;
wire  signed [31:0] sext_ln856_31_fu_25275_p1;
wire   [0:0] xor_ln896_68_fu_25403_p2;
wire   [0:0] xor_ln888_65_fu_25413_p2;
wire   [0:0] or_ln888_34_fu_25418_p2;
wire   [0:0] tmp_201_fu_25428_p3;
wire   [0:0] xor_ln890_32_fu_25436_p2;
wire   [0:0] or_ln890_34_fu_25442_p2;
wire   [0:0] carry_66_fu_25408_p2;
wire   [0:0] deleted_zeros_31_fu_25423_p2;
wire   [0:0] xor_ln895_68_fu_25458_p2;
wire   [0:0] or_ln895_34_fu_25464_p2;
wire   [0:0] xor_ln895_69_fu_25469_p2;
wire   [0:0] deleted_ones_34_fu_25448_p2;
wire   [0:0] xor_ln896_69_fu_25480_p2;
wire   [0:0] and_ln891_34_fu_25453_p2;
wire   [0:0] or_ln896_34_fu_25486_p2;
wire   [0:0] xor_ln896_277_fu_25492_p2;
wire   [0:0] overflow_34_fu_25474_p2;
wire   [0:0] underflow_34_fu_25498_p2;
wire   [0:0] or_ln346_34_fu_25511_p2;
wire   [31:0] select_ln346_68_fu_25503_p3;
wire  signed [31:0] sext_ln856_32_fu_25400_p1;
wire   [0:0] xor_ln896_70_fu_25525_p2;
wire   [0:0] xor_ln888_67_fu_25535_p2;
wire   [0:0] or_ln888_35_fu_25540_p2;
wire   [0:0] tmp_207_fu_25550_p3;
wire   [0:0] xor_ln890_33_fu_25558_p2;
wire   [0:0] or_ln890_35_fu_25564_p2;
wire   [0:0] carry_68_fu_25530_p2;
wire   [0:0] deleted_zeros_32_fu_25545_p2;
wire   [0:0] xor_ln895_70_fu_25580_p2;
wire   [0:0] or_ln895_35_fu_25586_p2;
wire   [0:0] xor_ln895_71_fu_25591_p2;
wire   [0:0] deleted_ones_35_fu_25570_p2;
wire   [0:0] xor_ln896_71_fu_25602_p2;
wire   [0:0] and_ln891_35_fu_25575_p2;
wire   [0:0] or_ln896_35_fu_25608_p2;
wire   [0:0] xor_ln896_278_fu_25614_p2;
wire   [0:0] overflow_35_fu_25596_p2;
wire   [0:0] underflow_35_fu_25620_p2;
wire   [0:0] or_ln346_35_fu_25633_p2;
wire   [31:0] select_ln346_70_fu_25625_p3;
wire   [27:0] zext_ln377_36_fu_25649_p1;
wire  signed [27:0] sext_ln823_33_fu_25646_p1;
wire  signed [27:0] p_Val2_107_fu_25652_p2;
wire   [0:0] p_Result_108_fu_25662_p3;
wire   [0:0] xor_ln896_72_fu_25670_p2;
wire   [0:0] xor_ln888_69_fu_25681_p2;
wire   [0:0] or_ln888_36_fu_25686_p2;
wire   [0:0] tmp_213_fu_25697_p3;
wire   [0:0] xor_ln890_34_fu_25705_p2;
wire   [0:0] or_ln890_36_fu_25711_p2;
wire   [0:0] carry_70_fu_25676_p2;
wire   [0:0] deleted_zeros_33_fu_25692_p2;
wire   [0:0] xor_ln895_72_fu_25727_p2;
wire   [0:0] or_ln895_36_fu_25733_p2;
wire   [0:0] xor_ln895_73_fu_25739_p2;
wire   [0:0] deleted_ones_36_fu_25717_p2;
wire   [0:0] xor_ln896_73_fu_25750_p2;
wire   [0:0] and_ln891_36_fu_25722_p2;
wire   [0:0] or_ln896_36_fu_25756_p2;
wire   [0:0] xor_ln896_279_fu_25762_p2;
wire   [0:0] overflow_36_fu_25744_p2;
wire   [0:0] underflow_36_fu_25768_p2;
wire   [0:0] or_ln346_36_fu_25781_p2;
wire   [31:0] select_ln346_72_fu_25773_p3;
wire  signed [31:0] sext_ln856_33_fu_25658_p1;
wire   [20:0] zext_ln377_37_fu_25798_p1;
wire  signed [20:0] sext_ln823_34_fu_25795_p1;
wire  signed [20:0] p_Val2_110_fu_25801_p2;
wire   [0:0] p_Result_111_fu_25811_p3;
wire   [0:0] xor_ln896_74_fu_25819_p2;
wire   [0:0] xor_ln888_71_fu_25830_p2;
wire   [0:0] or_ln888_37_fu_25835_p2;
wire   [0:0] tmp_219_fu_25846_p3;
wire   [0:0] xor_ln890_35_fu_25854_p2;
wire   [0:0] or_ln890_37_fu_25860_p2;
wire   [0:0] carry_72_fu_25825_p2;
wire   [0:0] deleted_zeros_34_fu_25841_p2;
wire   [0:0] xor_ln895_74_fu_25876_p2;
wire   [0:0] or_ln895_37_fu_25882_p2;
wire   [0:0] xor_ln895_75_fu_25888_p2;
wire   [0:0] deleted_ones_37_fu_25866_p2;
wire   [0:0] xor_ln896_75_fu_25899_p2;
wire   [0:0] and_ln891_37_fu_25871_p2;
wire   [0:0] or_ln896_37_fu_25905_p2;
wire   [0:0] xor_ln896_280_fu_25911_p2;
wire   [0:0] overflow_37_fu_25893_p2;
wire   [0:0] underflow_37_fu_25917_p2;
wire   [0:0] or_ln346_37_fu_25930_p2;
wire   [31:0] select_ln346_74_fu_25922_p3;
wire  signed [31:0] sext_ln856_34_fu_25807_p1;
wire   [18:0] zext_ln377_38_fu_25947_p1;
wire  signed [18:0] sext_ln823_35_fu_25944_p1;
wire  signed [18:0] p_Val2_113_fu_25950_p2;
wire   [0:0] p_Result_114_fu_25960_p3;
wire   [0:0] xor_ln896_76_fu_25968_p2;
wire   [0:0] xor_ln888_73_fu_25979_p2;
wire   [0:0] or_ln888_38_fu_25984_p2;
wire   [0:0] tmp_225_fu_25995_p3;
wire   [0:0] xor_ln890_36_fu_26003_p2;
wire   [0:0] or_ln890_38_fu_26009_p2;
wire   [0:0] carry_74_fu_25974_p2;
wire   [0:0] deleted_zeros_35_fu_25990_p2;
wire   [0:0] xor_ln895_76_fu_26025_p2;
wire   [0:0] or_ln895_38_fu_26031_p2;
wire   [0:0] xor_ln895_77_fu_26037_p2;
wire   [0:0] deleted_ones_38_fu_26015_p2;
wire   [0:0] xor_ln896_77_fu_26048_p2;
wire   [0:0] and_ln891_38_fu_26020_p2;
wire   [0:0] or_ln896_38_fu_26054_p2;
wire   [0:0] xor_ln896_281_fu_26060_p2;
wire   [0:0] overflow_38_fu_26042_p2;
wire   [0:0] underflow_38_fu_26066_p2;
wire   [0:0] or_ln346_38_fu_26079_p2;
wire   [31:0] select_ln346_76_fu_26071_p3;
wire  signed [31:0] sext_ln856_35_fu_25956_p1;
wire   [31:0] select_ln346_78_fu_26096_p3;
wire  signed [31:0] sext_ln856_36_fu_26093_p1;
wire   [19:0] zext_ln377_40_fu_26113_p1;
wire  signed [19:0] sext_ln823_37_fu_26110_p1;
wire  signed [19:0] p_Val2_119_fu_26116_p2;
wire   [0:0] p_Result_120_fu_26126_p3;
wire   [0:0] xor_ln896_80_fu_26134_p2;
wire   [0:0] xor_ln888_77_fu_26145_p2;
wire   [0:0] or_ln888_40_fu_26150_p2;
wire   [0:0] tmp_237_fu_26161_p3;
wire   [0:0] xor_ln890_38_fu_26169_p2;
wire   [0:0] or_ln890_40_fu_26175_p2;
wire   [0:0] carry_78_fu_26140_p2;
wire   [0:0] deleted_zeros_37_fu_26156_p2;
wire   [0:0] xor_ln895_80_fu_26191_p2;
wire   [0:0] or_ln895_40_fu_26197_p2;
wire   [0:0] xor_ln895_81_fu_26203_p2;
wire   [0:0] deleted_ones_40_fu_26181_p2;
wire   [0:0] xor_ln896_81_fu_26214_p2;
wire   [0:0] and_ln891_40_fu_26186_p2;
wire   [0:0] or_ln896_40_fu_26220_p2;
wire   [0:0] xor_ln896_283_fu_26226_p2;
wire   [0:0] overflow_40_fu_26208_p2;
wire   [0:0] underflow_40_fu_26232_p2;
wire   [0:0] or_ln346_40_fu_26245_p2;
wire   [31:0] select_ln346_80_fu_26237_p3;
wire  signed [31:0] sext_ln856_37_fu_26122_p1;
wire   [20:0] zext_ln377_41_fu_26262_p1;
wire  signed [20:0] sext_ln823_38_fu_26259_p1;
wire  signed [20:0] p_Val2_122_fu_26265_p2;
wire   [0:0] p_Result_123_fu_26275_p3;
wire   [0:0] xor_ln896_82_fu_26283_p2;
wire   [0:0] xor_ln888_79_fu_26294_p2;
wire   [0:0] or_ln888_41_fu_26299_p2;
wire   [0:0] tmp_243_fu_26310_p3;
wire   [0:0] xor_ln890_39_fu_26318_p2;
wire   [0:0] or_ln890_41_fu_26324_p2;
wire   [0:0] carry_80_fu_26289_p2;
wire   [0:0] deleted_zeros_38_fu_26305_p2;
wire   [0:0] xor_ln895_82_fu_26340_p2;
wire   [0:0] or_ln895_41_fu_26346_p2;
wire   [0:0] xor_ln895_83_fu_26352_p2;
wire   [0:0] deleted_ones_41_fu_26330_p2;
wire   [0:0] xor_ln896_83_fu_26363_p2;
wire   [0:0] and_ln891_41_fu_26335_p2;
wire   [0:0] or_ln896_41_fu_26369_p2;
wire   [0:0] xor_ln896_284_fu_26375_p2;
wire   [0:0] overflow_41_fu_26357_p2;
wire   [0:0] underflow_41_fu_26381_p2;
wire   [0:0] or_ln346_41_fu_26394_p2;
wire   [31:0] select_ln346_82_fu_26386_p3;
wire  signed [31:0] sext_ln856_38_fu_26271_p1;
wire   [19:0] zext_ln377_42_fu_26411_p1;
wire  signed [19:0] sext_ln823_39_fu_26408_p1;
wire  signed [19:0] p_Val2_125_fu_26414_p2;
wire   [0:0] p_Result_126_fu_26424_p3;
wire   [0:0] xor_ln896_84_fu_26432_p2;
wire   [0:0] xor_ln888_81_fu_26443_p2;
wire   [0:0] or_ln888_42_fu_26448_p2;
wire   [0:0] tmp_249_fu_26459_p3;
wire   [0:0] xor_ln890_40_fu_26467_p2;
wire   [0:0] or_ln890_42_fu_26473_p2;
wire   [0:0] carry_82_fu_26438_p2;
wire   [0:0] deleted_zeros_39_fu_26454_p2;
wire   [0:0] xor_ln895_84_fu_26489_p2;
wire   [0:0] or_ln895_42_fu_26495_p2;
wire   [0:0] xor_ln895_85_fu_26501_p2;
wire   [0:0] deleted_ones_42_fu_26479_p2;
wire   [0:0] xor_ln896_85_fu_26512_p2;
wire   [0:0] and_ln891_42_fu_26484_p2;
wire   [0:0] or_ln896_42_fu_26518_p2;
wire   [0:0] xor_ln896_285_fu_26524_p2;
wire   [0:0] overflow_42_fu_26506_p2;
wire   [0:0] underflow_42_fu_26530_p2;
wire   [0:0] or_ln346_42_fu_26543_p2;
wire   [31:0] select_ln346_84_fu_26535_p3;
wire  signed [31:0] sext_ln856_39_fu_26420_p1;
wire   [21:0] zext_ln377_43_fu_26560_p1;
wire  signed [21:0] sext_ln823_40_fu_26557_p1;
wire  signed [21:0] p_Val2_128_fu_26563_p2;
wire   [0:0] p_Result_129_fu_26573_p3;
wire   [0:0] xor_ln896_86_fu_26581_p2;
wire   [0:0] xor_ln888_83_fu_26592_p2;
wire   [0:0] or_ln888_43_fu_26597_p2;
wire   [0:0] tmp_255_fu_26608_p3;
wire   [0:0] xor_ln890_41_fu_26616_p2;
wire   [0:0] or_ln890_43_fu_26622_p2;
wire   [0:0] carry_84_fu_26587_p2;
wire   [0:0] deleted_zeros_40_fu_26603_p2;
wire   [0:0] xor_ln895_86_fu_26638_p2;
wire   [0:0] or_ln895_43_fu_26644_p2;
wire   [0:0] xor_ln895_87_fu_26650_p2;
wire   [0:0] deleted_ones_43_fu_26628_p2;
wire   [0:0] xor_ln896_87_fu_26661_p2;
wire   [0:0] and_ln891_43_fu_26633_p2;
wire   [0:0] or_ln896_43_fu_26667_p2;
wire   [0:0] xor_ln896_286_fu_26673_p2;
wire   [0:0] overflow_43_fu_26655_p2;
wire   [0:0] underflow_43_fu_26679_p2;
wire   [0:0] or_ln346_43_fu_26692_p2;
wire   [31:0] select_ln346_86_fu_26684_p3;
wire  signed [31:0] sext_ln856_40_fu_26569_p1;
wire   [29:0] zext_ln377_44_fu_26709_p1;
wire  signed [29:0] sext_ln823_41_fu_26706_p1;
wire  signed [29:0] p_Val2_131_fu_26712_p2;
wire   [0:0] p_Result_132_fu_26722_p3;
wire   [0:0] xor_ln896_88_fu_26730_p2;
wire   [0:0] xor_ln888_85_fu_26741_p2;
wire   [0:0] or_ln888_44_fu_26746_p2;
wire   [0:0] tmp_261_fu_26757_p3;
wire   [0:0] xor_ln890_42_fu_26765_p2;
wire   [0:0] or_ln890_44_fu_26771_p2;
wire   [0:0] carry_86_fu_26736_p2;
wire   [0:0] deleted_zeros_41_fu_26752_p2;
wire   [0:0] xor_ln895_88_fu_26787_p2;
wire   [0:0] or_ln895_44_fu_26793_p2;
wire   [0:0] xor_ln895_89_fu_26799_p2;
wire   [0:0] deleted_ones_44_fu_26777_p2;
wire   [0:0] xor_ln896_89_fu_26810_p2;
wire   [0:0] and_ln891_44_fu_26782_p2;
wire   [0:0] or_ln896_44_fu_26816_p2;
wire   [0:0] xor_ln896_287_fu_26822_p2;
wire   [0:0] overflow_44_fu_26804_p2;
wire   [0:0] underflow_44_fu_26828_p2;
wire   [0:0] or_ln346_44_fu_26841_p2;
wire   [31:0] select_ln346_88_fu_26833_p3;
wire  signed [31:0] sext_ln856_41_fu_26718_p1;
wire   [36:0] shl_ln1273_4_fu_26876_p3;
wire  signed [37:0] sext_ln70_30_fu_26873_p1;
wire  signed [37:0] sext_ln1273_4_fu_26883_p1;
wire   [37:0] r_V_42_fu_26887_p2;
wire   [13:0] p_Val2_133_fu_26901_p4;
wire   [14:0] zext_ln377_45_fu_26923_p1;
wire  signed [14:0] sext_ln823_42_fu_26911_p1;
wire   [0:0] p_Result_135_fu_26932_p3;
wire   [0:0] p_Result_134_fu_26915_p3;
wire   [0:0] xor_ln896_90_fu_26940_p2;
wire   [0:0] xor_ln888_87_fu_26960_p2;
wire   [0:0] Range2_all_ones_43_fu_26952_p3;
wire   [0:0] or_ln888_45_fu_26966_p2;
wire   [0:0] tmp_267_fu_26978_p3;
wire   [0:0] xor_ln890_43_fu_26986_p2;
wire   [0:0] or_ln890_45_fu_26992_p2;
wire   [0:0] carry_88_fu_26946_p2;
wire   [0:0] deleted_zeros_42_fu_26972_p2;
wire   [0:0] xor_ln895_90_fu_27010_p2;
wire   [0:0] p_Result_133_fu_26893_p3;
wire   [0:0] or_ln895_45_fu_27016_p2;
wire   [0:0] xor_ln895_91_fu_27022_p2;
wire   [0:0] deleted_ones_45_fu_26998_p2;
wire   [0:0] xor_ln896_91_fu_27034_p2;
wire   [0:0] and_ln891_45_fu_27004_p2;
wire   [0:0] or_ln896_45_fu_27040_p2;
wire   [0:0] xor_ln896_288_fu_27046_p2;
wire   [0:0] underflow_45_fu_27052_p2;
wire   [18:0] p_Val2_136_fu_27072_p4;
wire   [0:0] tmp_270_fu_27094_p3;
wire   [19:0] zext_ln377_46_fu_27102_p1;
wire  signed [19:0] sext_ln823_43_fu_27082_p1;
wire   [17:0] p_Val2_139_fu_27136_p4;
wire   [0:0] tmp_276_fu_27158_p3;
wire   [18:0] zext_ln377_47_fu_27166_p1;
wire  signed [18:0] sext_ln823_44_fu_27146_p1;
wire   [20:0] p_Val2_142_fu_27200_p4;
wire   [0:0] tmp_282_fu_27222_p3;
wire   [21:0] zext_ln377_48_fu_27230_p1;
wire  signed [21:0] sext_ln823_45_fu_27210_p1;
wire   [19:0] p_Val2_145_fu_27264_p4;
wire   [0:0] tmp_288_fu_27286_p3;
wire   [20:0] zext_ln377_49_fu_27294_p1;
wire  signed [20:0] sext_ln823_46_fu_27274_p1;
wire   [18:0] p_Val2_148_fu_27328_p4;
wire   [0:0] tmp_294_fu_27350_p3;
wire   [19:0] zext_ln377_50_fu_27358_p1;
wire  signed [19:0] sext_ln823_47_fu_27338_p1;
wire   [40:0] shl_ln1273_5_fu_27384_p3;
wire  signed [41:0] sext_ln1273_5_fu_27391_p1;
wire   [33:0] shl_ln1273_6_fu_27401_p3;
wire   [41:0] sub_ln1273_fu_27395_p2;
wire  signed [41:0] sext_ln1273_6_fu_27408_p1;
wire   [41:0] r_V_48_fu_27412_p2;
wire   [17:0] p_Val2_151_fu_27426_p4;
wire   [0:0] tmp_300_fu_27448_p3;
wire   [18:0] zext_ln377_51_fu_27456_p1;
wire  signed [18:0] sext_ln823_48_fu_27436_p1;
wire   [0:0] p_Result_153_fu_27466_p3;
wire   [0:0] p_Result_152_fu_27440_p3;
wire   [0:0] xor_ln896_102_fu_27474_p2;
wire   [0:0] xor_ln888_99_fu_27494_p2;
wire   [0:0] Range2_all_ones_49_fu_27486_p3;
wire   [0:0] or_ln888_51_fu_27500_p2;
wire   [0:0] tmp_303_fu_27512_p3;
wire   [0:0] xor_ln890_49_fu_27520_p2;
wire   [0:0] or_ln890_51_fu_27526_p2;
wire   [0:0] carry_100_fu_27480_p2;
wire   [0:0] deleted_zeros_48_fu_27506_p2;
wire   [0:0] xor_ln895_102_fu_27544_p2;
wire   [0:0] p_Result_151_fu_27418_p3;
wire   [0:0] or_ln895_51_fu_27550_p2;
wire   [0:0] xor_ln895_103_fu_27556_p2;
wire   [0:0] deleted_ones_51_fu_27532_p2;
wire   [0:0] xor_ln896_103_fu_27568_p2;
wire   [0:0] and_ln891_51_fu_27538_p2;
wire   [0:0] or_ln896_51_fu_27574_p2;
wire   [0:0] xor_ln896_294_fu_27580_p2;
wire   [0:0] underflow_51_fu_27586_p2;
wire   [18:0] p_Val2_154_fu_27606_p4;
wire   [0:0] tmp_306_fu_27628_p3;
wire   [19:0] zext_ln377_52_fu_27636_p1;
wire  signed [19:0] sext_ln823_49_fu_27616_p1;
wire   [32:0] shl_ln1273_7_fu_27662_p3;
wire  signed [41:0] sext_ln1273_7_fu_27669_p1;
wire   [41:0] r_V_50_fu_27673_p2;
wire   [17:0] p_Val2_157_fu_27687_p4;
wire   [0:0] tmp_312_fu_27709_p3;
wire   [18:0] zext_ln377_53_fu_27717_p1;
wire  signed [18:0] sext_ln823_50_fu_27697_p1;
wire   [0:0] p_Result_159_fu_27727_p3;
wire   [0:0] p_Result_158_fu_27701_p3;
wire   [0:0] xor_ln896_106_fu_27735_p2;
wire   [0:0] xor_ln888_103_fu_27755_p2;
wire   [0:0] Range2_all_ones_51_fu_27747_p3;
wire   [0:0] or_ln888_53_fu_27761_p2;
wire   [0:0] tmp_315_fu_27773_p3;
wire   [0:0] xor_ln890_51_fu_27781_p2;
wire   [0:0] or_ln890_53_fu_27787_p2;
wire   [0:0] carry_104_fu_27741_p2;
wire   [0:0] deleted_zeros_50_fu_27767_p2;
wire   [0:0] xor_ln895_106_fu_27805_p2;
wire   [0:0] p_Result_157_fu_27679_p3;
wire   [0:0] or_ln895_53_fu_27811_p2;
wire   [0:0] xor_ln895_107_fu_27817_p2;
wire   [0:0] deleted_ones_53_fu_27793_p2;
wire   [0:0] xor_ln896_107_fu_27829_p2;
wire   [0:0] and_ln891_53_fu_27799_p2;
wire   [0:0] or_ln896_53_fu_27835_p2;
wire   [0:0] xor_ln896_296_fu_27841_p2;
wire   [0:0] underflow_53_fu_27847_p2;
wire   [40:0] shl_ln1273_8_fu_28173_p3;
wire   [34:0] shl_ln1273_9_fu_28184_p3;
wire  signed [41:0] sext_ln1273_8_fu_28180_p1;
wire  signed [41:0] sext_ln1273_9_fu_28191_p1;
wire   [41:0] r_V_58_fu_28195_p2;
wire   [17:0] p_Val2_181_fu_28209_p4;
wire   [0:0] tmp_360_fu_28231_p3;
wire   [18:0] zext_ln377_61_fu_28239_p1;
wire  signed [18:0] sext_ln823_58_fu_28219_p1;
wire   [0:0] p_Result_183_fu_28249_p3;
wire   [0:0] p_Result_182_fu_28223_p3;
wire   [0:0] xor_ln896_122_fu_28257_p2;
wire   [0:0] xor_ln888_119_fu_28277_p2;
wire   [0:0] Range2_all_ones_59_fu_28269_p3;
wire   [0:0] or_ln888_61_fu_28283_p2;
wire   [0:0] tmp_363_fu_28295_p3;
wire   [0:0] xor_ln890_59_fu_28303_p2;
wire   [0:0] or_ln890_61_fu_28309_p2;
wire   [0:0] carry_120_fu_28263_p2;
wire   [0:0] deleted_zeros_58_fu_28289_p2;
wire   [0:0] xor_ln895_122_fu_28327_p2;
wire   [0:0] p_Result_181_fu_28201_p3;
wire   [0:0] or_ln895_61_fu_28333_p2;
wire   [0:0] xor_ln895_123_fu_28339_p2;
wire   [0:0] deleted_ones_61_fu_28315_p2;
wire   [0:0] xor_ln896_123_fu_28351_p2;
wire   [0:0] and_ln891_61_fu_28321_p2;
wire   [0:0] or_ln896_61_fu_28357_p2;
wire   [0:0] xor_ln896_304_fu_28363_p2;
wire   [0:0] underflow_61_fu_28369_p2;
wire  signed [31:0] rhs_18_fu_24420_p3;
wire  signed [32:0] sext_ln813_28_fu_28426_p1;
wire  signed [32:0] sext_ln813_27_fu_28423_p1;
wire   [32:0] ret_V_18_fu_28430_p2;
wire   [31:0] p_Val2_277_fu_28444_p2;
wire   [0:0] p_Result_277_fu_28436_p3;
wire   [0:0] p_Result_278_fu_28449_p3;
wire   [0:0] xor_ln895_180_fu_28457_p2;
wire   [0:0] xor_ln896_180_fu_28469_p2;
wire   [0:0] xor_ln302_36_fu_28481_p2;
wire   [0:0] overflow_99_fu_28463_p2;
wire   [0:0] xor_ln302_37_fu_28487_p2;
wire   [0:0] underflow_99_fu_28475_p2;
wire   [0:0] or_ln302_18_fu_28493_p2;
wire   [31:0] select_ln302_36_fu_28499_p3;
wire   [31:0] select_ln350_18_fu_28507_p3;
wire  signed [31:0] rhs_19_fu_24437_p3;
wire  signed [32:0] sext_ln813_30_fu_28526_p1;
wire  signed [32:0] sext_ln813_29_fu_28523_p1;
wire   [32:0] ret_V_19_fu_28530_p2;
wire   [31:0] p_Val2_279_fu_28544_p2;
wire   [0:0] p_Result_279_fu_28536_p3;
wire   [0:0] p_Result_280_fu_28549_p3;
wire   [0:0] xor_ln895_181_fu_28557_p2;
wire   [0:0] xor_ln896_181_fu_28569_p2;
wire   [0:0] xor_ln302_38_fu_28581_p2;
wire   [0:0] overflow_100_fu_28563_p2;
wire   [0:0] xor_ln302_39_fu_28587_p2;
wire   [0:0] underflow_100_fu_28575_p2;
wire   [0:0] or_ln302_19_fu_28593_p2;
wire   [31:0] select_ln302_38_fu_28599_p3;
wire   [31:0] select_ln350_19_fu_28607_p3;
wire   [0:0] xor_ln895_182_fu_28623_p2;
wire   [0:0] xor_ln896_182_fu_28633_p2;
wire   [0:0] xor_ln302_40_fu_28643_p2;
wire   [0:0] overflow_101_fu_28628_p2;
wire   [0:0] xor_ln302_41_fu_28647_p2;
wire   [0:0] underflow_101_fu_28638_p2;
wire   [0:0] or_ln302_20_fu_28653_p2;
wire   [31:0] select_ln302_40_fu_28659_p3;
wire   [31:0] select_ln350_20_fu_28666_p3;
wire  signed [31:0] rhs_21_fu_24454_p3;
wire  signed [32:0] sext_ln813_34_fu_28684_p1;
wire  signed [32:0] sext_ln813_33_fu_28681_p1;
wire   [32:0] ret_V_21_fu_28688_p2;
wire   [31:0] p_Val2_283_fu_28702_p2;
wire   [0:0] p_Result_283_fu_28694_p3;
wire   [0:0] p_Result_284_fu_28707_p3;
wire   [0:0] xor_ln895_183_fu_28715_p2;
wire   [0:0] xor_ln896_183_fu_28727_p2;
wire   [0:0] xor_ln302_42_fu_28739_p2;
wire   [0:0] overflow_102_fu_28721_p2;
wire   [0:0] xor_ln302_43_fu_28745_p2;
wire   [0:0] underflow_102_fu_28733_p2;
wire   [0:0] or_ln302_21_fu_28751_p2;
wire   [31:0] select_ln302_42_fu_28757_p3;
wire   [31:0] select_ln350_21_fu_28765_p3;
wire  signed [31:0] rhs_22_fu_24471_p3;
wire  signed [32:0] sext_ln813_36_fu_28784_p1;
wire  signed [32:0] sext_ln813_35_fu_28781_p1;
wire   [32:0] ret_V_22_fu_28788_p2;
wire   [31:0] p_Val2_285_fu_28802_p2;
wire   [0:0] p_Result_285_fu_28794_p3;
wire   [0:0] p_Result_286_fu_28807_p3;
wire   [0:0] xor_ln895_184_fu_28815_p2;
wire   [0:0] xor_ln896_184_fu_28827_p2;
wire   [0:0] xor_ln302_44_fu_28839_p2;
wire   [0:0] overflow_103_fu_28821_p2;
wire   [0:0] xor_ln302_45_fu_28845_p2;
wire   [0:0] underflow_103_fu_28833_p2;
wire   [0:0] or_ln302_22_fu_28851_p2;
wire   [31:0] select_ln302_44_fu_28857_p3;
wire   [31:0] select_ln350_22_fu_28865_p3;
wire  signed [31:0] rhs_23_fu_24488_p3;
wire  signed [32:0] sext_ln813_38_fu_28884_p1;
wire  signed [32:0] sext_ln813_37_fu_28881_p1;
wire   [32:0] ret_V_23_fu_28888_p2;
wire   [31:0] p_Val2_287_fu_28902_p2;
wire   [0:0] p_Result_287_fu_28894_p3;
wire   [0:0] p_Result_288_fu_28907_p3;
wire   [0:0] xor_ln895_185_fu_28915_p2;
wire   [0:0] xor_ln896_185_fu_28927_p2;
wire   [0:0] xor_ln302_46_fu_28939_p2;
wire   [0:0] overflow_104_fu_28921_p2;
wire   [0:0] xor_ln302_47_fu_28945_p2;
wire   [0:0] underflow_104_fu_28933_p2;
wire   [0:0] or_ln302_23_fu_28951_p2;
wire   [31:0] select_ln302_46_fu_28957_p3;
wire   [31:0] select_ln350_23_fu_28965_p3;
wire   [0:0] xor_ln895_186_fu_28981_p2;
wire   [0:0] xor_ln896_186_fu_28991_p2;
wire   [0:0] xor_ln302_48_fu_29001_p2;
wire   [0:0] overflow_105_fu_28986_p2;
wire   [0:0] xor_ln302_49_fu_29005_p2;
wire   [0:0] underflow_105_fu_28996_p2;
wire   [0:0] or_ln302_24_fu_29011_p2;
wire   [31:0] select_ln302_48_fu_29017_p3;
wire   [31:0] select_ln350_24_fu_29024_p3;
wire  signed [31:0] rhs_25_fu_24505_p3;
wire  signed [32:0] sext_ln813_42_fu_29042_p1;
wire  signed [32:0] sext_ln813_41_fu_29039_p1;
wire   [32:0] ret_V_25_fu_29046_p2;
wire   [31:0] p_Val2_291_fu_29060_p2;
wire   [0:0] p_Result_291_fu_29052_p3;
wire   [0:0] p_Result_292_fu_29065_p3;
wire   [0:0] xor_ln895_187_fu_29073_p2;
wire   [0:0] xor_ln896_187_fu_29085_p2;
wire   [0:0] xor_ln302_50_fu_29097_p2;
wire   [0:0] overflow_106_fu_29079_p2;
wire   [0:0] xor_ln302_51_fu_29103_p2;
wire   [0:0] underflow_106_fu_29091_p2;
wire   [0:0] or_ln302_25_fu_29109_p2;
wire   [31:0] select_ln302_50_fu_29115_p3;
wire   [31:0] select_ln350_25_fu_29123_p3;
wire  signed [31:0] rhs_26_fu_24522_p3;
wire  signed [32:0] sext_ln813_44_fu_29142_p1;
wire  signed [32:0] sext_ln813_43_fu_29139_p1;
wire   [32:0] ret_V_26_fu_29146_p2;
wire   [31:0] p_Val2_293_fu_29160_p2;
wire   [0:0] p_Result_293_fu_29152_p3;
wire   [0:0] p_Result_294_fu_29165_p3;
wire   [0:0] xor_ln895_188_fu_29173_p2;
wire   [0:0] xor_ln896_188_fu_29185_p2;
wire   [0:0] xor_ln302_52_fu_29197_p2;
wire   [0:0] overflow_107_fu_29179_p2;
wire   [0:0] xor_ln302_53_fu_29203_p2;
wire   [0:0] underflow_107_fu_29191_p2;
wire   [0:0] or_ln302_26_fu_29209_p2;
wire   [31:0] select_ln302_52_fu_29215_p3;
wire   [31:0] select_ln350_26_fu_29223_p3;
wire  signed [31:0] lhs_18_fu_28515_p3;
wire  signed [31:0] rhs_27_fu_24643_p3;
wire  signed [32:0] sext_ln813_46_fu_29243_p1;
wire  signed [32:0] sext_ln813_45_fu_29239_p1;
wire   [32:0] ret_V_27_fu_29247_p2;
wire   [31:0] p_Val2_295_fu_29261_p2;
wire   [0:0] p_Result_295_fu_29253_p3;
wire   [0:0] p_Result_296_fu_29267_p3;
wire   [0:0] xor_ln895_189_fu_29275_p2;
wire   [0:0] xor_ln896_189_fu_29287_p2;
wire   [0:0] xor_ln302_54_fu_29299_p2;
wire   [0:0] overflow_108_fu_29281_p2;
wire   [0:0] xor_ln302_55_fu_29305_p2;
wire   [0:0] underflow_108_fu_29293_p2;
wire   [0:0] or_ln302_27_fu_29311_p2;
wire   [31:0] select_ln302_54_fu_29317_p3;
wire   [31:0] select_ln350_27_fu_29325_p3;
wire  signed [31:0] lhs_19_fu_28615_p3;
wire  signed [31:0] rhs_28_fu_24767_p3;
wire  signed [32:0] sext_ln813_48_fu_29345_p1;
wire  signed [32:0] sext_ln813_47_fu_29341_p1;
wire   [32:0] ret_V_28_fu_29349_p2;
wire   [31:0] p_Val2_297_fu_29363_p2;
wire   [0:0] p_Result_297_fu_29355_p3;
wire   [0:0] p_Result_298_fu_29369_p3;
wire   [0:0] xor_ln895_190_fu_29377_p2;
wire   [0:0] xor_ln896_190_fu_29389_p2;
wire   [0:0] xor_ln302_56_fu_29401_p2;
wire   [0:0] overflow_109_fu_29383_p2;
wire   [0:0] xor_ln302_57_fu_29407_p2;
wire   [0:0] underflow_109_fu_29395_p2;
wire   [0:0] or_ln302_28_fu_29413_p2;
wire   [31:0] select_ln302_56_fu_29419_p3;
wire   [31:0] select_ln350_28_fu_29427_p3;
wire  signed [31:0] lhs_20_fu_28673_p3;
wire  signed [31:0] rhs_29_fu_24892_p3;
wire  signed [32:0] sext_ln813_50_fu_29447_p1;
wire  signed [32:0] sext_ln813_49_fu_29443_p1;
wire   [32:0] ret_V_29_fu_29451_p2;
wire   [31:0] p_Val2_299_fu_29465_p2;
wire   [0:0] p_Result_299_fu_29457_p3;
wire   [0:0] p_Result_300_fu_29471_p3;
wire   [0:0] xor_ln895_191_fu_29479_p2;
wire   [0:0] xor_ln896_191_fu_29491_p2;
wire   [0:0] xor_ln302_58_fu_29503_p2;
wire   [0:0] overflow_110_fu_29485_p2;
wire   [0:0] xor_ln302_59_fu_29509_p2;
wire   [0:0] underflow_110_fu_29497_p2;
wire   [0:0] or_ln302_29_fu_29515_p2;
wire   [31:0] select_ln302_58_fu_29521_p3;
wire   [31:0] select_ln350_29_fu_29529_p3;
wire  signed [31:0] lhs_21_fu_28773_p3;
wire  signed [31:0] rhs_30_fu_25017_p3;
wire  signed [32:0] sext_ln813_52_fu_29549_p1;
wire  signed [32:0] sext_ln813_51_fu_29545_p1;
wire   [32:0] ret_V_30_fu_29553_p2;
wire   [31:0] p_Val2_301_fu_29567_p2;
wire   [0:0] p_Result_301_fu_29559_p3;
wire   [0:0] p_Result_302_fu_29573_p3;
wire   [0:0] xor_ln895_192_fu_29581_p2;
wire   [0:0] xor_ln896_192_fu_29593_p2;
wire   [0:0] xor_ln302_60_fu_29605_p2;
wire   [0:0] overflow_111_fu_29587_p2;
wire   [0:0] xor_ln302_61_fu_29611_p2;
wire   [0:0] underflow_111_fu_29599_p2;
wire   [0:0] or_ln302_30_fu_29617_p2;
wire   [31:0] select_ln302_60_fu_29623_p3;
wire   [31:0] select_ln350_30_fu_29631_p3;
wire  signed [31:0] lhs_22_fu_28873_p3;
wire  signed [31:0] rhs_31_fu_25142_p3;
wire  signed [32:0] sext_ln813_54_fu_29651_p1;
wire  signed [32:0] sext_ln813_53_fu_29647_p1;
wire   [32:0] ret_V_31_fu_29655_p2;
wire   [31:0] p_Val2_303_fu_29669_p2;
wire   [0:0] p_Result_303_fu_29661_p3;
wire   [0:0] p_Result_304_fu_29675_p3;
wire   [0:0] xor_ln895_193_fu_29683_p2;
wire   [0:0] xor_ln896_193_fu_29695_p2;
wire   [0:0] xor_ln302_62_fu_29707_p2;
wire   [0:0] overflow_112_fu_29689_p2;
wire   [0:0] xor_ln302_63_fu_29713_p2;
wire   [0:0] underflow_112_fu_29701_p2;
wire   [0:0] or_ln302_31_fu_29719_p2;
wire   [31:0] select_ln302_62_fu_29725_p3;
wire   [31:0] select_ln350_31_fu_29733_p3;
wire  signed [31:0] lhs_23_fu_28973_p3;
wire  signed [31:0] rhs_32_fu_25267_p3;
wire  signed [32:0] sext_ln813_56_fu_29753_p1;
wire  signed [32:0] sext_ln813_55_fu_29749_p1;
wire   [32:0] ret_V_32_fu_29757_p2;
wire   [31:0] p_Val2_305_fu_29771_p2;
wire   [0:0] p_Result_305_fu_29763_p3;
wire   [0:0] p_Result_306_fu_29777_p3;
wire   [0:0] xor_ln895_194_fu_29785_p2;
wire   [0:0] xor_ln896_194_fu_29797_p2;
wire   [0:0] xor_ln302_64_fu_29809_p2;
wire   [0:0] overflow_113_fu_29791_p2;
wire   [0:0] xor_ln302_65_fu_29815_p2;
wire   [0:0] underflow_113_fu_29803_p2;
wire   [0:0] or_ln302_32_fu_29821_p2;
wire   [31:0] select_ln302_64_fu_29827_p3;
wire   [31:0] select_ln350_32_fu_29835_p3;
wire  signed [31:0] lhs_24_fu_29031_p3;
wire  signed [31:0] rhs_33_fu_25392_p3;
wire  signed [32:0] sext_ln813_58_fu_29855_p1;
wire  signed [32:0] sext_ln813_57_fu_29851_p1;
wire   [32:0] ret_V_33_fu_29859_p2;
wire   [31:0] p_Val2_307_fu_29873_p2;
wire   [0:0] p_Result_307_fu_29865_p3;
wire   [0:0] p_Result_308_fu_29879_p3;
wire   [0:0] xor_ln895_195_fu_29887_p2;
wire   [0:0] xor_ln896_195_fu_29899_p2;
wire   [0:0] xor_ln302_66_fu_29911_p2;
wire   [0:0] overflow_114_fu_29893_p2;
wire   [0:0] xor_ln302_67_fu_29917_p2;
wire   [0:0] underflow_114_fu_29905_p2;
wire   [0:0] or_ln302_33_fu_29923_p2;
wire   [31:0] select_ln302_66_fu_29929_p3;
wire   [31:0] select_ln350_33_fu_29937_p3;
wire  signed [31:0] lhs_25_fu_29131_p3;
wire  signed [31:0] rhs_34_fu_25517_p3;
wire  signed [32:0] sext_ln813_60_fu_29957_p1;
wire  signed [32:0] sext_ln813_59_fu_29953_p1;
wire   [32:0] ret_V_34_fu_29961_p2;
wire   [31:0] p_Val2_309_fu_29975_p2;
wire   [0:0] p_Result_309_fu_29967_p3;
wire   [0:0] p_Result_310_fu_29981_p3;
wire   [0:0] xor_ln895_196_fu_29989_p2;
wire   [0:0] xor_ln896_196_fu_30001_p2;
wire   [0:0] xor_ln302_68_fu_30013_p2;
wire   [0:0] overflow_115_fu_29995_p2;
wire   [0:0] xor_ln302_69_fu_30019_p2;
wire   [0:0] underflow_115_fu_30007_p2;
wire   [0:0] or_ln302_34_fu_30025_p2;
wire   [31:0] select_ln302_68_fu_30031_p3;
wire   [31:0] select_ln350_34_fu_30039_p3;
wire  signed [31:0] lhs_26_fu_29231_p3;
wire  signed [31:0] rhs_35_fu_25639_p3;
wire  signed [32:0] sext_ln813_62_fu_30059_p1;
wire  signed [32:0] sext_ln813_61_fu_30055_p1;
wire   [32:0] ret_V_35_fu_30063_p2;
wire   [31:0] p_Val2_311_fu_30077_p2;
wire   [0:0] p_Result_311_fu_30069_p3;
wire   [0:0] p_Result_312_fu_30083_p3;
wire   [0:0] xor_ln895_197_fu_30091_p2;
wire   [0:0] xor_ln896_197_fu_30103_p2;
wire   [0:0] xor_ln302_70_fu_30115_p2;
wire   [0:0] overflow_116_fu_30097_p2;
wire   [0:0] xor_ln302_71_fu_30121_p2;
wire   [0:0] underflow_116_fu_30109_p2;
wire   [0:0] or_ln302_35_fu_30127_p2;
wire   [31:0] select_ln302_70_fu_30133_p3;
wire   [31:0] select_ln350_35_fu_30141_p3;
wire  signed [31:0] lhs_27_fu_29333_p3;
wire  signed [31:0] rhs_36_fu_25787_p3;
wire  signed [32:0] sext_ln813_64_fu_30161_p1;
wire  signed [32:0] sext_ln813_63_fu_30157_p1;
wire   [32:0] ret_V_36_fu_30165_p2;
wire  signed [31:0] lhs_28_fu_29435_p3;
wire  signed [31:0] rhs_37_fu_25936_p3;
wire  signed [32:0] sext_ln813_66_fu_30197_p1;
wire  signed [32:0] sext_ln813_65_fu_30193_p1;
wire   [32:0] ret_V_37_fu_30201_p2;
wire  signed [31:0] lhs_29_fu_29537_p3;
wire  signed [31:0] rhs_38_fu_26085_p3;
wire  signed [32:0] sext_ln813_68_fu_30233_p1;
wire  signed [32:0] sext_ln813_67_fu_30229_p1;
wire   [32:0] ret_V_38_fu_30237_p2;
wire   [31:0] p_Val2_317_fu_30251_p2;
wire   [0:0] p_Result_317_fu_30243_p3;
wire   [0:0] p_Result_318_fu_30257_p3;
wire   [0:0] xor_ln895_200_fu_30265_p2;
wire   [0:0] xor_ln896_200_fu_30277_p2;
wire   [0:0] xor_ln302_76_fu_30289_p2;
wire   [0:0] overflow_119_fu_30271_p2;
wire   [0:0] xor_ln302_77_fu_30295_p2;
wire   [0:0] underflow_119_fu_30283_p2;
wire   [0:0] or_ln302_38_fu_30301_p2;
wire   [31:0] select_ln302_76_fu_30307_p3;
wire   [31:0] select_ln350_38_fu_30315_p3;
wire  signed [31:0] lhs_30_fu_29639_p3;
wire  signed [31:0] rhs_39_fu_26103_p3;
wire  signed [32:0] sext_ln813_70_fu_30335_p1;
wire  signed [32:0] sext_ln813_69_fu_30331_p1;
wire   [32:0] ret_V_39_fu_30339_p2;
wire  signed [31:0] lhs_31_fu_29741_p3;
wire  signed [31:0] rhs_40_fu_26251_p3;
wire  signed [32:0] sext_ln813_72_fu_30371_p1;
wire  signed [32:0] sext_ln813_71_fu_30367_p1;
wire   [32:0] ret_V_40_fu_30375_p2;
wire  signed [31:0] lhs_32_fu_29843_p3;
wire  signed [31:0] rhs_41_fu_26400_p3;
wire  signed [32:0] sext_ln813_74_fu_30407_p1;
wire  signed [32:0] sext_ln813_73_fu_30403_p1;
wire   [32:0] ret_V_41_fu_30411_p2;
wire  signed [31:0] lhs_33_fu_29945_p3;
wire  signed [31:0] rhs_42_fu_26549_p3;
wire  signed [32:0] sext_ln813_76_fu_30443_p1;
wire  signed [32:0] sext_ln813_75_fu_30439_p1;
wire   [32:0] ret_V_42_fu_30447_p2;
wire   [31:0] p_Val2_325_fu_30461_p2;
wire   [0:0] p_Result_325_fu_30453_p3;
wire   [0:0] p_Result_326_fu_30467_p3;
wire   [0:0] xor_ln895_204_fu_30475_p2;
wire   [0:0] xor_ln896_204_fu_30487_p2;
wire   [0:0] xor_ln302_84_fu_30499_p2;
wire   [0:0] overflow_123_fu_30481_p2;
wire   [0:0] xor_ln302_85_fu_30505_p2;
wire   [0:0] underflow_123_fu_30493_p2;
wire   [0:0] or_ln302_42_fu_30511_p2;
wire   [31:0] select_ln302_84_fu_30517_p3;
wire   [31:0] select_ln350_42_fu_30525_p3;
wire  signed [31:0] lhs_34_fu_30047_p3;
wire  signed [31:0] rhs_43_fu_26698_p3;
wire  signed [32:0] sext_ln813_78_fu_30545_p1;
wire  signed [32:0] sext_ln813_77_fu_30541_p1;
wire   [32:0] ret_V_43_fu_30549_p2;
wire  signed [31:0] lhs_35_fu_30149_p3;
wire  signed [31:0] rhs_44_fu_26847_p3;
wire  signed [32:0] sext_ln813_80_fu_30581_p1;
wire  signed [32:0] sext_ln813_79_fu_30577_p1;
wire   [32:0] ret_V_44_fu_30585_p2;
wire   [31:0] select_ln346_90_fu_30616_p3;
wire  signed [31:0] sext_ln856_42_fu_30613_p1;
wire   [0:0] xor_ln896_92_fu_30633_p2;
wire   [0:0] xor_ln888_89_fu_30643_p2;
wire   [0:0] or_ln888_46_fu_30648_p2;
wire   [0:0] tmp_273_fu_30658_p3;
wire   [0:0] xor_ln890_44_fu_30666_p2;
wire   [0:0] or_ln890_46_fu_30672_p2;
wire   [0:0] carry_90_fu_30638_p2;
wire   [0:0] deleted_zeros_43_fu_30653_p2;
wire   [0:0] xor_ln895_92_fu_30688_p2;
wire   [0:0] or_ln895_46_fu_30694_p2;
wire   [0:0] xor_ln895_93_fu_30699_p2;
wire   [0:0] deleted_ones_46_fu_30678_p2;
wire   [0:0] xor_ln896_93_fu_30710_p2;
wire   [0:0] and_ln891_46_fu_30683_p2;
wire   [0:0] or_ln896_46_fu_30716_p2;
wire   [0:0] xor_ln896_289_fu_30722_p2;
wire   [0:0] overflow_46_fu_30704_p2;
wire   [0:0] underflow_46_fu_30728_p2;
wire   [0:0] or_ln346_46_fu_30741_p2;
wire   [31:0] select_ln346_92_fu_30733_p3;
wire  signed [31:0] sext_ln856_43_fu_30630_p1;
wire   [0:0] xor_ln896_94_fu_30758_p2;
wire   [0:0] xor_ln888_91_fu_30768_p2;
wire   [0:0] or_ln888_47_fu_30773_p2;
wire   [0:0] tmp_279_fu_30783_p3;
wire   [0:0] xor_ln890_45_fu_30791_p2;
wire   [0:0] or_ln890_47_fu_30797_p2;
wire   [0:0] carry_92_fu_30763_p2;
wire   [0:0] deleted_zeros_44_fu_30778_p2;
wire   [0:0] xor_ln895_94_fu_30813_p2;
wire   [0:0] or_ln895_47_fu_30819_p2;
wire   [0:0] xor_ln895_95_fu_30824_p2;
wire   [0:0] deleted_ones_47_fu_30803_p2;
wire   [0:0] xor_ln896_95_fu_30835_p2;
wire   [0:0] and_ln891_47_fu_30808_p2;
wire   [0:0] or_ln896_47_fu_30841_p2;
wire   [0:0] xor_ln896_290_fu_30847_p2;
wire   [0:0] overflow_47_fu_30829_p2;
wire   [0:0] underflow_47_fu_30853_p2;
wire   [0:0] or_ln346_47_fu_30866_p2;
wire   [31:0] select_ln346_94_fu_30858_p3;
wire  signed [31:0] sext_ln856_44_fu_30755_p1;
wire   [0:0] xor_ln896_96_fu_30883_p2;
wire   [0:0] xor_ln888_93_fu_30893_p2;
wire   [0:0] or_ln888_48_fu_30898_p2;
wire   [0:0] tmp_285_fu_30908_p3;
wire   [0:0] xor_ln890_46_fu_30916_p2;
wire   [0:0] or_ln890_48_fu_30922_p2;
wire   [0:0] carry_94_fu_30888_p2;
wire   [0:0] deleted_zeros_45_fu_30903_p2;
wire   [0:0] xor_ln895_96_fu_30938_p2;
wire   [0:0] or_ln895_48_fu_30944_p2;
wire   [0:0] xor_ln895_97_fu_30949_p2;
wire   [0:0] deleted_ones_48_fu_30928_p2;
wire   [0:0] xor_ln896_97_fu_30960_p2;
wire   [0:0] and_ln891_48_fu_30933_p2;
wire   [0:0] or_ln896_48_fu_30966_p2;
wire   [0:0] xor_ln896_291_fu_30972_p2;
wire   [0:0] overflow_48_fu_30954_p2;
wire   [0:0] underflow_48_fu_30978_p2;
wire   [0:0] or_ln346_48_fu_30991_p2;
wire   [31:0] select_ln346_96_fu_30983_p3;
wire  signed [31:0] sext_ln856_45_fu_30880_p1;
wire   [0:0] xor_ln896_98_fu_31008_p2;
wire   [0:0] xor_ln888_95_fu_31018_p2;
wire   [0:0] or_ln888_49_fu_31023_p2;
wire   [0:0] tmp_291_fu_31033_p3;
wire   [0:0] xor_ln890_47_fu_31041_p2;
wire   [0:0] or_ln890_49_fu_31047_p2;
wire   [0:0] carry_96_fu_31013_p2;
wire   [0:0] deleted_zeros_46_fu_31028_p2;
wire   [0:0] xor_ln895_98_fu_31063_p2;
wire   [0:0] or_ln895_49_fu_31069_p2;
wire   [0:0] xor_ln895_99_fu_31074_p2;
wire   [0:0] deleted_ones_49_fu_31053_p2;
wire   [0:0] xor_ln896_99_fu_31085_p2;
wire   [0:0] and_ln891_49_fu_31058_p2;
wire   [0:0] or_ln896_49_fu_31091_p2;
wire   [0:0] xor_ln896_292_fu_31097_p2;
wire   [0:0] overflow_49_fu_31079_p2;
wire   [0:0] underflow_49_fu_31103_p2;
wire   [0:0] or_ln346_49_fu_31116_p2;
wire   [31:0] select_ln346_98_fu_31108_p3;
wire  signed [31:0] sext_ln856_46_fu_31005_p1;
wire   [0:0] xor_ln896_100_fu_31133_p2;
wire   [0:0] xor_ln888_97_fu_31143_p2;
wire   [0:0] or_ln888_50_fu_31148_p2;
wire   [0:0] tmp_297_fu_31158_p3;
wire   [0:0] xor_ln890_48_fu_31166_p2;
wire   [0:0] or_ln890_50_fu_31172_p2;
wire   [0:0] carry_98_fu_31138_p2;
wire   [0:0] deleted_zeros_47_fu_31153_p2;
wire   [0:0] xor_ln895_100_fu_31188_p2;
wire   [0:0] or_ln895_50_fu_31194_p2;
wire   [0:0] xor_ln895_101_fu_31199_p2;
wire   [0:0] deleted_ones_50_fu_31178_p2;
wire   [0:0] xor_ln896_101_fu_31210_p2;
wire   [0:0] and_ln891_50_fu_31183_p2;
wire   [0:0] or_ln896_50_fu_31216_p2;
wire   [0:0] xor_ln896_293_fu_31222_p2;
wire   [0:0] overflow_50_fu_31204_p2;
wire   [0:0] underflow_50_fu_31228_p2;
wire   [0:0] or_ln346_50_fu_31241_p2;
wire   [31:0] select_ln346_100_fu_31233_p3;
wire  signed [31:0] sext_ln856_47_fu_31130_p1;
wire   [31:0] select_ln346_102_fu_31258_p3;
wire  signed [31:0] sext_ln856_48_fu_31255_p1;
wire   [0:0] xor_ln896_104_fu_31275_p2;
wire   [0:0] xor_ln888_101_fu_31285_p2;
wire   [0:0] or_ln888_52_fu_31290_p2;
wire   [0:0] tmp_309_fu_31300_p3;
wire   [0:0] xor_ln890_50_fu_31308_p2;
wire   [0:0] or_ln890_52_fu_31314_p2;
wire   [0:0] carry_102_fu_31280_p2;
wire   [0:0] deleted_zeros_49_fu_31295_p2;
wire   [0:0] xor_ln895_104_fu_31330_p2;
wire   [0:0] or_ln895_52_fu_31336_p2;
wire   [0:0] xor_ln895_105_fu_31341_p2;
wire   [0:0] deleted_ones_52_fu_31320_p2;
wire   [0:0] xor_ln896_105_fu_31352_p2;
wire   [0:0] and_ln891_52_fu_31325_p2;
wire   [0:0] or_ln896_52_fu_31358_p2;
wire   [0:0] xor_ln896_295_fu_31364_p2;
wire   [0:0] overflow_52_fu_31346_p2;
wire   [0:0] underflow_52_fu_31370_p2;
wire   [0:0] or_ln346_52_fu_31383_p2;
wire   [31:0] select_ln346_104_fu_31375_p3;
wire  signed [31:0] sext_ln856_49_fu_31272_p1;
wire   [31:0] select_ln346_106_fu_31400_p3;
wire  signed [31:0] sext_ln856_50_fu_31397_p1;
wire   [19:0] zext_ln377_54_fu_31417_p1;
wire  signed [19:0] sext_ln823_51_fu_31414_p1;
wire  signed [19:0] p_Val2_161_fu_31420_p2;
wire   [0:0] p_Result_162_fu_31430_p3;
wire   [0:0] xor_ln896_108_fu_31438_p2;
wire   [0:0] xor_ln888_105_fu_31449_p2;
wire   [0:0] or_ln888_54_fu_31454_p2;
wire   [0:0] tmp_321_fu_31465_p3;
wire   [0:0] xor_ln890_52_fu_31473_p2;
wire   [0:0] or_ln890_54_fu_31479_p2;
wire   [0:0] carry_106_fu_31444_p2;
wire   [0:0] deleted_zeros_51_fu_31460_p2;
wire   [0:0] xor_ln895_108_fu_31495_p2;
wire   [0:0] or_ln895_54_fu_31501_p2;
wire   [0:0] xor_ln895_109_fu_31507_p2;
wire   [0:0] deleted_ones_54_fu_31485_p2;
wire   [0:0] xor_ln896_109_fu_31518_p2;
wire   [0:0] and_ln891_54_fu_31490_p2;
wire   [0:0] or_ln896_54_fu_31524_p2;
wire   [0:0] xor_ln896_297_fu_31530_p2;
wire   [0:0] overflow_54_fu_31512_p2;
wire   [0:0] underflow_54_fu_31536_p2;
wire   [0:0] or_ln346_54_fu_31549_p2;
wire   [31:0] select_ln346_108_fu_31541_p3;
wire  signed [31:0] sext_ln856_51_fu_31426_p1;
wire   [18:0] zext_ln377_55_fu_31566_p1;
wire  signed [18:0] sext_ln823_52_fu_31563_p1;
wire  signed [18:0] p_Val2_164_fu_31569_p2;
wire   [0:0] p_Result_165_fu_31579_p3;
wire   [0:0] xor_ln896_110_fu_31587_p2;
wire   [0:0] xor_ln888_107_fu_31598_p2;
wire   [0:0] or_ln888_55_fu_31603_p2;
wire   [0:0] tmp_327_fu_31614_p3;
wire   [0:0] xor_ln890_53_fu_31622_p2;
wire   [0:0] or_ln890_55_fu_31628_p2;
wire   [0:0] carry_108_fu_31593_p2;
wire   [0:0] deleted_zeros_52_fu_31609_p2;
wire   [0:0] xor_ln895_110_fu_31644_p2;
wire   [0:0] or_ln895_55_fu_31650_p2;
wire   [0:0] xor_ln895_111_fu_31656_p2;
wire   [0:0] deleted_ones_55_fu_31634_p2;
wire   [0:0] xor_ln896_111_fu_31667_p2;
wire   [0:0] and_ln891_55_fu_31639_p2;
wire   [0:0] or_ln896_55_fu_31673_p2;
wire   [0:0] xor_ln896_298_fu_31679_p2;
wire   [0:0] overflow_55_fu_31661_p2;
wire   [0:0] underflow_55_fu_31685_p2;
wire   [0:0] or_ln346_55_fu_31698_p2;
wire   [31:0] select_ln346_110_fu_31690_p3;
wire  signed [31:0] sext_ln856_52_fu_31575_p1;
wire   [20:0] zext_ln377_56_fu_31715_p1;
wire  signed [20:0] sext_ln823_53_fu_31712_p1;
wire  signed [20:0] p_Val2_167_fu_31718_p2;
wire   [0:0] p_Result_168_fu_31728_p3;
wire   [0:0] xor_ln896_112_fu_31736_p2;
wire   [0:0] xor_ln888_109_fu_31747_p2;
wire   [0:0] or_ln888_56_fu_31752_p2;
wire   [0:0] tmp_333_fu_31763_p3;
wire   [0:0] xor_ln890_54_fu_31771_p2;
wire   [0:0] or_ln890_56_fu_31777_p2;
wire   [0:0] carry_110_fu_31742_p2;
wire   [0:0] deleted_zeros_53_fu_31758_p2;
wire   [0:0] xor_ln895_112_fu_31793_p2;
wire   [0:0] or_ln895_56_fu_31799_p2;
wire   [0:0] xor_ln895_113_fu_31805_p2;
wire   [0:0] deleted_ones_56_fu_31783_p2;
wire   [0:0] xor_ln896_113_fu_31816_p2;
wire   [0:0] and_ln891_56_fu_31788_p2;
wire   [0:0] or_ln896_56_fu_31822_p2;
wire   [0:0] xor_ln896_299_fu_31828_p2;
wire   [0:0] overflow_56_fu_31810_p2;
wire   [0:0] underflow_56_fu_31834_p2;
wire   [0:0] or_ln346_56_fu_31847_p2;
wire   [31:0] select_ln346_112_fu_31839_p3;
wire  signed [31:0] sext_ln856_53_fu_31724_p1;
wire   [21:0] zext_ln377_57_fu_31864_p1;
wire  signed [21:0] sext_ln823_54_fu_31861_p1;
wire  signed [21:0] p_Val2_170_fu_31867_p2;
wire   [0:0] p_Result_171_fu_31877_p3;
wire   [0:0] xor_ln896_114_fu_31885_p2;
wire   [0:0] xor_ln888_111_fu_31896_p2;
wire   [0:0] or_ln888_57_fu_31901_p2;
wire   [0:0] tmp_339_fu_31912_p3;
wire   [0:0] xor_ln890_55_fu_31920_p2;
wire   [0:0] or_ln890_57_fu_31926_p2;
wire   [0:0] carry_112_fu_31891_p2;
wire   [0:0] deleted_zeros_54_fu_31907_p2;
wire   [0:0] xor_ln895_114_fu_31942_p2;
wire   [0:0] or_ln895_57_fu_31948_p2;
wire   [0:0] xor_ln895_115_fu_31954_p2;
wire   [0:0] deleted_ones_57_fu_31932_p2;
wire   [0:0] xor_ln896_115_fu_31965_p2;
wire   [0:0] and_ln891_57_fu_31937_p2;
wire   [0:0] or_ln896_57_fu_31971_p2;
wire   [0:0] xor_ln896_300_fu_31977_p2;
wire   [0:0] overflow_57_fu_31959_p2;
wire   [0:0] underflow_57_fu_31983_p2;
wire   [0:0] or_ln346_57_fu_31996_p2;
wire   [31:0] select_ln346_114_fu_31988_p3;
wire  signed [31:0] sext_ln856_54_fu_31873_p1;
wire   [21:0] zext_ln377_58_fu_32013_p1;
wire  signed [21:0] sext_ln823_55_fu_32010_p1;
wire  signed [21:0] p_Val2_173_fu_32016_p2;
wire   [0:0] p_Result_174_fu_32026_p3;
wire   [0:0] xor_ln896_116_fu_32034_p2;
wire   [0:0] xor_ln888_113_fu_32045_p2;
wire   [0:0] or_ln888_58_fu_32050_p2;
wire   [0:0] tmp_345_fu_32061_p3;
wire   [0:0] xor_ln890_56_fu_32069_p2;
wire   [0:0] or_ln890_58_fu_32075_p2;
wire   [0:0] carry_114_fu_32040_p2;
wire   [0:0] deleted_zeros_55_fu_32056_p2;
wire   [0:0] xor_ln895_116_fu_32091_p2;
wire   [0:0] or_ln895_58_fu_32097_p2;
wire   [0:0] xor_ln895_117_fu_32103_p2;
wire   [0:0] deleted_ones_58_fu_32081_p2;
wire   [0:0] xor_ln896_117_fu_32114_p2;
wire   [0:0] and_ln891_58_fu_32086_p2;
wire   [0:0] or_ln896_58_fu_32120_p2;
wire   [0:0] xor_ln896_301_fu_32126_p2;
wire   [0:0] overflow_58_fu_32108_p2;
wire   [0:0] underflow_58_fu_32132_p2;
wire   [0:0] or_ln346_58_fu_32145_p2;
wire   [31:0] select_ln346_116_fu_32137_p3;
wire  signed [31:0] sext_ln856_55_fu_32022_p1;
wire   [20:0] zext_ln377_59_fu_32162_p1;
wire  signed [20:0] sext_ln823_56_fu_32159_p1;
wire  signed [20:0] p_Val2_176_fu_32165_p2;
wire   [0:0] p_Result_177_fu_32175_p3;
wire   [0:0] xor_ln896_118_fu_32183_p2;
wire   [0:0] xor_ln888_115_fu_32194_p2;
wire   [0:0] or_ln888_59_fu_32199_p2;
wire   [0:0] tmp_351_fu_32210_p3;
wire   [0:0] xor_ln890_57_fu_32218_p2;
wire   [0:0] or_ln890_59_fu_32224_p2;
wire   [0:0] carry_116_fu_32189_p2;
wire   [0:0] deleted_zeros_56_fu_32205_p2;
wire   [0:0] xor_ln895_118_fu_32240_p2;
wire   [0:0] or_ln895_59_fu_32246_p2;
wire   [0:0] xor_ln895_119_fu_32252_p2;
wire   [0:0] deleted_ones_59_fu_32230_p2;
wire   [0:0] xor_ln896_119_fu_32263_p2;
wire   [0:0] and_ln891_59_fu_32235_p2;
wire   [0:0] or_ln896_59_fu_32269_p2;
wire   [0:0] xor_ln896_302_fu_32275_p2;
wire   [0:0] overflow_59_fu_32257_p2;
wire   [0:0] underflow_59_fu_32281_p2;
wire   [0:0] or_ln346_59_fu_32294_p2;
wire   [31:0] select_ln346_118_fu_32286_p3;
wire  signed [31:0] sext_ln856_56_fu_32171_p1;
wire   [21:0] zext_ln377_60_fu_32311_p1;
wire  signed [21:0] sext_ln823_57_fu_32308_p1;
wire  signed [21:0] p_Val2_179_fu_32314_p2;
wire   [0:0] p_Result_180_fu_32324_p3;
wire   [0:0] xor_ln896_120_fu_32332_p2;
wire   [0:0] xor_ln888_117_fu_32343_p2;
wire   [0:0] or_ln888_60_fu_32348_p2;
wire   [0:0] tmp_357_fu_32359_p3;
wire   [0:0] xor_ln890_58_fu_32367_p2;
wire   [0:0] or_ln890_60_fu_32373_p2;
wire   [0:0] carry_118_fu_32338_p2;
wire   [0:0] deleted_zeros_57_fu_32354_p2;
wire   [0:0] xor_ln895_120_fu_32389_p2;
wire   [0:0] or_ln895_60_fu_32395_p2;
wire   [0:0] xor_ln895_121_fu_32401_p2;
wire   [0:0] deleted_ones_60_fu_32379_p2;
wire   [0:0] xor_ln896_121_fu_32412_p2;
wire   [0:0] and_ln891_60_fu_32384_p2;
wire   [0:0] or_ln896_60_fu_32418_p2;
wire   [0:0] xor_ln896_303_fu_32424_p2;
wire   [0:0] overflow_60_fu_32406_p2;
wire   [0:0] underflow_60_fu_32430_p2;
wire   [0:0] or_ln346_60_fu_32443_p2;
wire   [31:0] select_ln346_120_fu_32435_p3;
wire  signed [31:0] sext_ln856_57_fu_32320_p1;
wire   [31:0] select_ln346_122_fu_32460_p3;
wire  signed [31:0] sext_ln856_58_fu_32457_p1;
wire   [20:0] zext_ln377_62_fu_32477_p1;
wire  signed [20:0] sext_ln823_59_fu_32474_p1;
wire  signed [20:0] p_Val2_185_fu_32480_p2;
wire   [0:0] p_Result_186_fu_32490_p3;
wire   [0:0] xor_ln896_124_fu_32498_p2;
wire   [0:0] xor_ln888_121_fu_32509_p2;
wire   [0:0] or_ln888_62_fu_32514_p2;
wire   [0:0] tmp_369_fu_32525_p3;
wire   [0:0] xor_ln890_60_fu_32533_p2;
wire   [0:0] or_ln890_62_fu_32539_p2;
wire   [0:0] carry_122_fu_32504_p2;
wire   [0:0] deleted_zeros_59_fu_32520_p2;
wire   [0:0] xor_ln895_124_fu_32555_p2;
wire   [0:0] or_ln895_62_fu_32561_p2;
wire   [0:0] xor_ln895_125_fu_32567_p2;
wire   [0:0] deleted_ones_62_fu_32545_p2;
wire   [0:0] xor_ln896_125_fu_32578_p2;
wire   [0:0] and_ln891_62_fu_32550_p2;
wire   [0:0] or_ln896_62_fu_32584_p2;
wire   [0:0] xor_ln896_305_fu_32590_p2;
wire   [0:0] overflow_62_fu_32572_p2;
wire   [0:0] underflow_62_fu_32596_p2;
wire   [0:0] or_ln346_62_fu_32609_p2;
wire   [31:0] select_ln346_124_fu_32601_p3;
wire  signed [31:0] sext_ln856_59_fu_32486_p1;
wire   [17:0] p_Val2_187_fu_32648_p4;
wire   [0:0] tmp_372_fu_32670_p3;
wire   [18:0] zext_ln377_63_fu_32678_p1;
wire  signed [18:0] sext_ln823_60_fu_32658_p1;
wire   [18:0] p_Val2_190_fu_32712_p4;
wire   [0:0] tmp_378_fu_32734_p3;
wire   [19:0] zext_ln377_64_fu_32742_p1;
wire  signed [19:0] sext_ln823_61_fu_32722_p1;
wire   [19:0] p_Val2_193_fu_32776_p4;
wire   [0:0] tmp_384_fu_32798_p3;
wire   [20:0] zext_ln377_65_fu_32806_p1;
wire  signed [20:0] sext_ln823_62_fu_32786_p1;
wire   [17:0] p_Val2_196_fu_32840_p4;
wire   [0:0] tmp_390_fu_32862_p3;
wire   [18:0] zext_ln377_66_fu_32870_p1;
wire  signed [18:0] sext_ln823_63_fu_32850_p1;
wire   [19:0] p_Val2_199_fu_32904_p4;
wire   [0:0] tmp_396_fu_32926_p3;
wire   [20:0] zext_ln377_67_fu_32934_p1;
wire  signed [20:0] sext_ln823_64_fu_32914_p1;
wire   [37:0] shl_ln1273_s_fu_32960_p3;
wire  signed [38:0] sext_ln1273_10_fu_32967_p1;
wire   [38:0] r_V_65_fu_32971_p2;
wire   [14:0] p_Val2_202_fu_32985_p4;
wire   [0:0] tmp_402_fu_33007_p3;
wire   [15:0] zext_ln377_68_fu_33015_p1;
wire  signed [15:0] sext_ln823_65_fu_32995_p1;
wire   [0:0] p_Result_204_fu_33025_p3;
wire   [0:0] p_Result_203_fu_32999_p3;
wire   [0:0] xor_ln896_136_fu_33033_p2;
wire   [0:0] xor_ln888_133_fu_33053_p2;
wire   [0:0] Range2_all_ones_66_fu_33045_p3;
wire   [0:0] or_ln888_68_fu_33059_p2;
wire   [0:0] tmp_405_fu_33071_p3;
wire   [0:0] xor_ln890_66_fu_33079_p2;
wire   [0:0] or_ln890_68_fu_33085_p2;
wire   [0:0] carry_134_fu_33039_p2;
wire   [0:0] deleted_zeros_65_fu_33065_p2;
wire   [0:0] xor_ln895_136_fu_33103_p2;
wire   [0:0] p_Result_202_fu_32977_p3;
wire   [0:0] or_ln895_68_fu_33109_p2;
wire   [0:0] xor_ln895_137_fu_33115_p2;
wire   [0:0] deleted_ones_68_fu_33091_p2;
wire   [0:0] xor_ln896_137_fu_33127_p2;
wire   [0:0] and_ln891_68_fu_33097_p2;
wire   [0:0] or_ln896_68_fu_33133_p2;
wire   [0:0] xor_ln896_311_fu_33139_p2;
wire   [0:0] underflow_68_fu_33145_p2;
wire   [18:0] p_Val2_205_fu_33165_p4;
wire   [0:0] tmp_408_fu_33187_p3;
wire   [19:0] zext_ln377_69_fu_33195_p1;
wire  signed [19:0] sext_ln823_66_fu_33175_p1;
wire   [19:0] p_Val2_208_fu_33229_p4;
wire   [0:0] tmp_414_fu_33251_p3;
wire   [20:0] zext_ln377_70_fu_33259_p1;
wire  signed [20:0] sext_ln823_67_fu_33239_p1;
wire   [17:0] p_Val2_211_fu_33293_p4;
wire   [0:0] tmp_420_fu_33315_p3;
wire   [18:0] zext_ln377_71_fu_33323_p1;
wire  signed [18:0] sext_ln823_68_fu_33303_p1;
wire   [38:0] shl_ln1273_10_fu_33546_p3;
wire   [35:0] shl_ln1273_11_fu_33557_p3;
wire  signed [39:0] sext_ln1273_11_fu_33553_p1;
wire  signed [39:0] sext_ln1273_12_fu_33564_p1;
wire   [39:0] r_V_73_fu_33568_p2;
wire   [15:0] p_Val2_226_fu_33582_p4;
wire   [0:0] tmp_450_fu_33604_p3;
wire   [16:0] zext_ln377_76_fu_33612_p1;
wire  signed [16:0] sext_ln823_73_fu_33592_p1;
wire   [0:0] p_Result_228_fu_33622_p3;
wire   [0:0] p_Result_227_fu_33596_p3;
wire   [0:0] xor_ln896_152_fu_33630_p2;
wire   [0:0] xor_ln888_149_fu_33650_p2;
wire   [0:0] Range2_all_ones_74_fu_33642_p3;
wire   [0:0] or_ln888_76_fu_33656_p2;
wire   [0:0] tmp_453_fu_33668_p3;
wire   [0:0] xor_ln890_74_fu_33676_p2;
wire   [0:0] or_ln890_76_fu_33682_p2;
wire   [0:0] carry_150_fu_33636_p2;
wire   [0:0] deleted_zeros_73_fu_33662_p2;
wire   [0:0] xor_ln895_152_fu_33700_p2;
wire   [0:0] p_Result_226_fu_33574_p3;
wire   [0:0] or_ln895_76_fu_33706_p2;
wire   [0:0] xor_ln895_153_fu_33712_p2;
wire   [0:0] deleted_ones_76_fu_33688_p2;
wire   [0:0] xor_ln896_153_fu_33724_p2;
wire   [0:0] and_ln891_76_fu_33694_p2;
wire   [0:0] or_ln896_76_fu_33730_p2;
wire   [0:0] xor_ln896_319_fu_33736_p2;
wire   [0:0] underflow_76_fu_33742_p2;
wire   [0:0] xor_ln895_198_fu_33922_p2;
wire   [0:0] xor_ln896_198_fu_33932_p2;
wire   [0:0] xor_ln302_72_fu_33942_p2;
wire   [0:0] overflow_117_fu_33927_p2;
wire   [0:0] xor_ln302_73_fu_33946_p2;
wire   [0:0] underflow_117_fu_33937_p2;
wire   [0:0] or_ln302_36_fu_33952_p2;
wire   [31:0] select_ln302_72_fu_33958_p3;
wire   [31:0] select_ln350_36_fu_33965_p3;
wire   [0:0] xor_ln895_199_fu_33980_p2;
wire   [0:0] xor_ln896_199_fu_33990_p2;
wire   [0:0] xor_ln302_74_fu_34000_p2;
wire   [0:0] overflow_118_fu_33985_p2;
wire   [0:0] xor_ln302_75_fu_34004_p2;
wire   [0:0] underflow_118_fu_33995_p2;
wire   [0:0] or_ln302_37_fu_34010_p2;
wire   [31:0] select_ln302_74_fu_34016_p3;
wire   [31:0] select_ln350_37_fu_34023_p3;
wire   [0:0] xor_ln895_201_fu_34038_p2;
wire   [0:0] xor_ln896_201_fu_34048_p2;
wire   [0:0] xor_ln302_78_fu_34058_p2;
wire   [0:0] overflow_120_fu_34043_p2;
wire   [0:0] xor_ln302_79_fu_34062_p2;
wire   [0:0] underflow_120_fu_34053_p2;
wire   [0:0] or_ln302_39_fu_34068_p2;
wire   [31:0] select_ln302_78_fu_34074_p3;
wire   [31:0] select_ln350_39_fu_34081_p3;
wire   [0:0] xor_ln895_202_fu_34096_p2;
wire   [0:0] xor_ln896_202_fu_34106_p2;
wire   [0:0] xor_ln302_80_fu_34116_p2;
wire   [0:0] overflow_121_fu_34101_p2;
wire   [0:0] xor_ln302_81_fu_34120_p2;
wire   [0:0] underflow_121_fu_34111_p2;
wire   [0:0] or_ln302_40_fu_34126_p2;
wire   [31:0] select_ln302_80_fu_34132_p3;
wire   [31:0] select_ln350_40_fu_34139_p3;
wire   [0:0] xor_ln895_203_fu_34154_p2;
wire   [0:0] xor_ln896_203_fu_34164_p2;
wire   [0:0] xor_ln302_82_fu_34174_p2;
wire   [0:0] overflow_122_fu_34159_p2;
wire   [0:0] xor_ln302_83_fu_34178_p2;
wire   [0:0] underflow_122_fu_34169_p2;
wire   [0:0] or_ln302_41_fu_34184_p2;
wire   [31:0] select_ln302_82_fu_34190_p3;
wire   [31:0] select_ln350_41_fu_34197_p3;
wire   [0:0] xor_ln895_205_fu_34212_p2;
wire   [0:0] xor_ln896_205_fu_34222_p2;
wire   [0:0] xor_ln302_86_fu_34232_p2;
wire   [0:0] overflow_124_fu_34217_p2;
wire   [0:0] xor_ln302_87_fu_34236_p2;
wire   [0:0] underflow_124_fu_34227_p2;
wire   [0:0] or_ln302_43_fu_34242_p2;
wire   [31:0] select_ln302_86_fu_34248_p3;
wire   [31:0] select_ln350_43_fu_34255_p3;
wire   [0:0] xor_ln895_206_fu_34270_p2;
wire   [0:0] xor_ln896_206_fu_34280_p2;
wire   [0:0] xor_ln302_88_fu_34290_p2;
wire   [0:0] overflow_125_fu_34275_p2;
wire   [0:0] xor_ln302_89_fu_34294_p2;
wire   [0:0] underflow_125_fu_34285_p2;
wire   [0:0] or_ln302_44_fu_34300_p2;
wire   [31:0] select_ln302_88_fu_34306_p3;
wire   [31:0] select_ln350_44_fu_34313_p3;
wire  signed [31:0] lhs_36_fu_33972_p3;
wire  signed [31:0] rhs_45_fu_30623_p3;
wire  signed [32:0] sext_ln813_82_fu_34332_p1;
wire  signed [32:0] sext_ln813_81_fu_34328_p1;
wire   [32:0] ret_V_45_fu_34336_p2;
wire   [31:0] p_Val2_331_fu_34350_p2;
wire   [0:0] p_Result_331_fu_34342_p3;
wire   [0:0] p_Result_332_fu_34356_p3;
wire   [0:0] xor_ln895_207_fu_34364_p2;
wire   [0:0] xor_ln896_207_fu_34376_p2;
wire   [0:0] xor_ln302_90_fu_34388_p2;
wire   [0:0] overflow_126_fu_34370_p2;
wire   [0:0] xor_ln302_91_fu_34394_p2;
wire   [0:0] underflow_126_fu_34382_p2;
wire   [0:0] or_ln302_45_fu_34400_p2;
wire   [31:0] select_ln302_90_fu_34406_p3;
wire   [31:0] select_ln350_45_fu_34414_p3;
wire  signed [31:0] lhs_37_fu_34030_p3;
wire  signed [31:0] rhs_46_fu_30747_p3;
wire  signed [32:0] sext_ln813_84_fu_34434_p1;
wire  signed [32:0] sext_ln813_83_fu_34430_p1;
wire   [32:0] ret_V_46_fu_34438_p2;
wire   [31:0] p_Val2_333_fu_34452_p2;
wire   [0:0] p_Result_333_fu_34444_p3;
wire   [0:0] p_Result_334_fu_34458_p3;
wire   [0:0] xor_ln895_208_fu_34466_p2;
wire   [0:0] xor_ln896_208_fu_34478_p2;
wire   [0:0] xor_ln302_92_fu_34490_p2;
wire   [0:0] overflow_127_fu_34472_p2;
wire   [0:0] xor_ln302_93_fu_34496_p2;
wire   [0:0] underflow_127_fu_34484_p2;
wire   [0:0] or_ln302_46_fu_34502_p2;
wire   [31:0] select_ln302_92_fu_34508_p3;
wire   [31:0] select_ln350_46_fu_34516_p3;
wire  signed [31:0] rhs_47_fu_30872_p3;
wire  signed [32:0] sext_ln813_86_fu_34535_p1;
wire  signed [32:0] sext_ln813_85_fu_34532_p1;
wire   [32:0] ret_V_47_fu_34539_p2;
wire   [31:0] p_Val2_335_fu_34553_p2;
wire   [0:0] p_Result_335_fu_34545_p3;
wire   [0:0] p_Result_336_fu_34558_p3;
wire   [0:0] xor_ln895_209_fu_34566_p2;
wire   [0:0] xor_ln896_209_fu_34578_p2;
wire   [0:0] xor_ln302_94_fu_34590_p2;
wire   [0:0] overflow_128_fu_34572_p2;
wire   [0:0] xor_ln302_95_fu_34596_p2;
wire   [0:0] underflow_128_fu_34584_p2;
wire   [0:0] or_ln302_47_fu_34602_p2;
wire   [31:0] select_ln302_94_fu_34608_p3;
wire   [31:0] select_ln350_47_fu_34616_p3;
wire  signed [31:0] lhs_39_fu_34088_p3;
wire  signed [31:0] rhs_48_fu_30997_p3;
wire  signed [32:0] sext_ln813_88_fu_34636_p1;
wire  signed [32:0] sext_ln813_87_fu_34632_p1;
wire   [32:0] ret_V_48_fu_34640_p2;
wire   [31:0] p_Val2_337_fu_34654_p2;
wire   [0:0] p_Result_337_fu_34646_p3;
wire   [0:0] p_Result_338_fu_34660_p3;
wire   [0:0] xor_ln895_210_fu_34668_p2;
wire   [0:0] xor_ln896_210_fu_34680_p2;
wire   [0:0] xor_ln302_96_fu_34692_p2;
wire   [0:0] overflow_129_fu_34674_p2;
wire   [0:0] xor_ln302_97_fu_34698_p2;
wire   [0:0] underflow_129_fu_34686_p2;
wire   [0:0] or_ln302_48_fu_34704_p2;
wire   [31:0] select_ln302_96_fu_34710_p3;
wire   [31:0] select_ln350_48_fu_34718_p3;
wire  signed [31:0] lhs_40_fu_34146_p3;
wire  signed [31:0] rhs_49_fu_31122_p3;
wire  signed [32:0] sext_ln813_90_fu_34738_p1;
wire  signed [32:0] sext_ln813_89_fu_34734_p1;
wire   [32:0] ret_V_49_fu_34742_p2;
wire   [31:0] p_Val2_339_fu_34756_p2;
wire   [0:0] p_Result_339_fu_34748_p3;
wire   [0:0] p_Result_340_fu_34762_p3;
wire   [0:0] xor_ln895_211_fu_34770_p2;
wire   [0:0] xor_ln896_211_fu_34782_p2;
wire   [0:0] xor_ln302_98_fu_34794_p2;
wire   [0:0] overflow_130_fu_34776_p2;
wire   [0:0] xor_ln302_99_fu_34800_p2;
wire   [0:0] underflow_130_fu_34788_p2;
wire   [0:0] or_ln302_49_fu_34806_p2;
wire   [31:0] select_ln302_98_fu_34812_p3;
wire   [31:0] select_ln350_49_fu_34820_p3;
wire  signed [31:0] lhs_41_fu_34204_p3;
wire  signed [31:0] rhs_50_fu_31247_p3;
wire  signed [32:0] sext_ln813_92_fu_34840_p1;
wire  signed [32:0] sext_ln813_91_fu_34836_p1;
wire   [32:0] ret_V_50_fu_34844_p2;
wire   [31:0] p_Val2_341_fu_34858_p2;
wire   [0:0] p_Result_341_fu_34850_p3;
wire   [0:0] p_Result_342_fu_34864_p3;
wire   [0:0] xor_ln895_212_fu_34872_p2;
wire   [0:0] xor_ln896_212_fu_34884_p2;
wire   [0:0] xor_ln302_100_fu_34896_p2;
wire   [0:0] overflow_131_fu_34878_p2;
wire   [0:0] xor_ln302_101_fu_34902_p2;
wire   [0:0] underflow_131_fu_34890_p2;
wire   [0:0] or_ln302_50_fu_34908_p2;
wire   [31:0] select_ln302_100_fu_34914_p3;
wire   [31:0] select_ln350_50_fu_34922_p3;
wire  signed [31:0] rhs_51_fu_31265_p3;
wire  signed [32:0] sext_ln813_94_fu_34941_p1;
wire  signed [32:0] sext_ln813_93_fu_34938_p1;
wire   [32:0] ret_V_51_fu_34945_p2;
wire   [31:0] p_Val2_343_fu_34959_p2;
wire   [0:0] p_Result_343_fu_34951_p3;
wire   [0:0] p_Result_344_fu_34964_p3;
wire   [0:0] xor_ln895_213_fu_34972_p2;
wire   [0:0] xor_ln896_213_fu_34984_p2;
wire   [0:0] xor_ln302_102_fu_34996_p2;
wire   [0:0] overflow_132_fu_34978_p2;
wire   [0:0] xor_ln302_103_fu_35002_p2;
wire   [0:0] underflow_132_fu_34990_p2;
wire   [0:0] or_ln302_51_fu_35008_p2;
wire   [31:0] select_ln302_102_fu_35014_p3;
wire   [31:0] select_ln350_51_fu_35022_p3;
wire  signed [31:0] lhs_43_fu_34262_p3;
wire  signed [31:0] rhs_52_fu_31389_p3;
wire  signed [32:0] sext_ln813_96_fu_35042_p1;
wire  signed [32:0] sext_ln813_95_fu_35038_p1;
wire   [32:0] ret_V_52_fu_35046_p2;
wire   [31:0] p_Val2_345_fu_35060_p2;
wire   [0:0] p_Result_345_fu_35052_p3;
wire   [0:0] p_Result_346_fu_35066_p3;
wire   [0:0] xor_ln895_214_fu_35074_p2;
wire   [0:0] xor_ln896_214_fu_35086_p2;
wire   [0:0] xor_ln302_104_fu_35098_p2;
wire   [0:0] overflow_133_fu_35080_p2;
wire   [0:0] xor_ln302_105_fu_35104_p2;
wire   [0:0] underflow_133_fu_35092_p2;
wire   [0:0] or_ln302_52_fu_35110_p2;
wire   [31:0] select_ln302_104_fu_35116_p3;
wire   [31:0] select_ln350_52_fu_35124_p3;
wire  signed [31:0] lhs_44_fu_34320_p3;
wire  signed [31:0] rhs_53_fu_31407_p3;
wire  signed [32:0] sext_ln813_98_fu_35144_p1;
wire  signed [32:0] sext_ln813_97_fu_35140_p1;
wire   [32:0] ret_V_53_fu_35148_p2;
wire   [31:0] p_Val2_347_fu_35162_p2;
wire   [0:0] p_Result_347_fu_35154_p3;
wire   [0:0] p_Result_348_fu_35168_p3;
wire   [0:0] xor_ln895_215_fu_35176_p2;
wire   [0:0] xor_ln896_215_fu_35188_p2;
wire   [0:0] xor_ln302_106_fu_35200_p2;
wire   [0:0] overflow_134_fu_35182_p2;
wire   [0:0] xor_ln302_107_fu_35206_p2;
wire   [0:0] underflow_134_fu_35194_p2;
wire   [0:0] or_ln302_53_fu_35212_p2;
wire   [31:0] select_ln302_106_fu_35218_p3;
wire   [31:0] select_ln350_53_fu_35226_p3;
wire  signed [31:0] lhs_45_fu_34422_p3;
wire  signed [31:0] rhs_54_fu_31555_p3;
wire  signed [32:0] sext_ln813_100_fu_35246_p1;
wire  signed [32:0] sext_ln813_99_fu_35242_p1;
wire   [32:0] ret_V_54_fu_35250_p2;
wire   [31:0] p_Val2_349_fu_35264_p2;
wire   [0:0] p_Result_349_fu_35256_p3;
wire   [0:0] p_Result_350_fu_35270_p3;
wire   [0:0] xor_ln895_216_fu_35278_p2;
wire   [0:0] xor_ln896_216_fu_35290_p2;
wire   [0:0] xor_ln302_108_fu_35302_p2;
wire   [0:0] overflow_135_fu_35284_p2;
wire   [0:0] xor_ln302_109_fu_35308_p2;
wire   [0:0] underflow_135_fu_35296_p2;
wire   [0:0] or_ln302_54_fu_35314_p2;
wire   [31:0] select_ln302_108_fu_35320_p3;
wire   [31:0] select_ln350_54_fu_35328_p3;
wire  signed [31:0] lhs_46_fu_34524_p3;
wire  signed [31:0] rhs_55_fu_31704_p3;
wire  signed [32:0] sext_ln813_102_fu_35348_p1;
wire  signed [32:0] sext_ln813_101_fu_35344_p1;
wire   [32:0] ret_V_55_fu_35352_p2;
wire   [31:0] p_Val2_351_fu_35366_p2;
wire   [0:0] p_Result_351_fu_35358_p3;
wire   [0:0] p_Result_352_fu_35372_p3;
wire   [0:0] xor_ln895_217_fu_35380_p2;
wire   [0:0] xor_ln896_217_fu_35392_p2;
wire   [0:0] xor_ln302_110_fu_35404_p2;
wire   [0:0] overflow_136_fu_35386_p2;
wire   [0:0] xor_ln302_111_fu_35410_p2;
wire   [0:0] underflow_136_fu_35398_p2;
wire   [0:0] or_ln302_55_fu_35416_p2;
wire   [31:0] select_ln302_110_fu_35422_p3;
wire   [31:0] select_ln350_55_fu_35430_p3;
wire  signed [31:0] lhs_47_fu_34624_p3;
wire  signed [31:0] rhs_56_fu_31853_p3;
wire  signed [32:0] sext_ln813_104_fu_35450_p1;
wire  signed [32:0] sext_ln813_103_fu_35446_p1;
wire   [32:0] ret_V_56_fu_35454_p2;
wire   [31:0] p_Val2_353_fu_35468_p2;
wire   [0:0] p_Result_353_fu_35460_p3;
wire   [0:0] p_Result_354_fu_35474_p3;
wire   [0:0] xor_ln895_218_fu_35482_p2;
wire   [0:0] xor_ln896_218_fu_35494_p2;
wire   [0:0] xor_ln302_112_fu_35506_p2;
wire   [0:0] overflow_137_fu_35488_p2;
wire   [0:0] xor_ln302_113_fu_35512_p2;
wire   [0:0] underflow_137_fu_35500_p2;
wire   [0:0] or_ln302_56_fu_35518_p2;
wire   [31:0] select_ln302_112_fu_35524_p3;
wire   [31:0] select_ln350_56_fu_35532_p3;
wire  signed [31:0] lhs_48_fu_34726_p3;
wire  signed [31:0] rhs_57_fu_32002_p3;
wire  signed [32:0] sext_ln813_106_fu_35552_p1;
wire  signed [32:0] sext_ln813_105_fu_35548_p1;
wire   [32:0] ret_V_57_fu_35556_p2;
wire   [31:0] p_Val2_355_fu_35570_p2;
wire   [0:0] p_Result_355_fu_35562_p3;
wire   [0:0] p_Result_356_fu_35576_p3;
wire   [0:0] xor_ln895_219_fu_35584_p2;
wire   [0:0] xor_ln896_219_fu_35596_p2;
wire   [0:0] xor_ln302_114_fu_35608_p2;
wire   [0:0] overflow_138_fu_35590_p2;
wire   [0:0] xor_ln302_115_fu_35614_p2;
wire   [0:0] underflow_138_fu_35602_p2;
wire   [0:0] or_ln302_57_fu_35620_p2;
wire   [31:0] select_ln302_114_fu_35626_p3;
wire   [31:0] select_ln350_57_fu_35634_p3;
wire  signed [31:0] lhs_49_fu_34828_p3;
wire  signed [31:0] rhs_58_fu_32151_p3;
wire  signed [32:0] sext_ln813_108_fu_35654_p1;
wire  signed [32:0] sext_ln813_107_fu_35650_p1;
wire   [32:0] ret_V_58_fu_35658_p2;
wire   [31:0] p_Val2_357_fu_35672_p2;
wire   [0:0] p_Result_357_fu_35664_p3;
wire   [0:0] p_Result_358_fu_35678_p3;
wire   [0:0] xor_ln895_220_fu_35686_p2;
wire   [0:0] xor_ln896_220_fu_35698_p2;
wire   [0:0] xor_ln302_116_fu_35710_p2;
wire   [0:0] overflow_139_fu_35692_p2;
wire   [0:0] xor_ln302_117_fu_35716_p2;
wire   [0:0] underflow_139_fu_35704_p2;
wire   [0:0] or_ln302_58_fu_35722_p2;
wire   [31:0] select_ln302_116_fu_35728_p3;
wire   [31:0] select_ln350_58_fu_35736_p3;
wire  signed [31:0] lhs_50_fu_34930_p3;
wire  signed [31:0] rhs_59_fu_32300_p3;
wire  signed [32:0] sext_ln813_110_fu_35756_p1;
wire  signed [32:0] sext_ln813_109_fu_35752_p1;
wire   [32:0] ret_V_59_fu_35760_p2;
wire   [31:0] p_Val2_359_fu_35774_p2;
wire   [0:0] p_Result_359_fu_35766_p3;
wire   [0:0] p_Result_360_fu_35780_p3;
wire   [0:0] xor_ln895_221_fu_35788_p2;
wire   [0:0] xor_ln896_221_fu_35800_p2;
wire   [0:0] xor_ln302_118_fu_35812_p2;
wire   [0:0] overflow_140_fu_35794_p2;
wire   [0:0] xor_ln302_119_fu_35818_p2;
wire   [0:0] underflow_140_fu_35806_p2;
wire   [0:0] or_ln302_59_fu_35824_p2;
wire   [31:0] select_ln302_118_fu_35830_p3;
wire   [31:0] select_ln350_59_fu_35838_p3;
wire  signed [31:0] lhs_51_fu_35030_p3;
wire  signed [31:0] rhs_60_fu_32449_p3;
wire  signed [32:0] sext_ln813_112_fu_35858_p1;
wire  signed [32:0] sext_ln813_111_fu_35854_p1;
wire   [32:0] ret_V_60_fu_35862_p2;
wire   [31:0] p_Val2_361_fu_35876_p2;
wire   [0:0] p_Result_361_fu_35868_p3;
wire   [0:0] p_Result_362_fu_35882_p3;
wire   [0:0] xor_ln895_222_fu_35890_p2;
wire   [0:0] xor_ln896_222_fu_35902_p2;
wire   [0:0] xor_ln302_120_fu_35914_p2;
wire   [0:0] overflow_141_fu_35896_p2;
wire   [0:0] xor_ln302_121_fu_35920_p2;
wire   [0:0] underflow_141_fu_35908_p2;
wire   [0:0] or_ln302_60_fu_35926_p2;
wire   [31:0] select_ln302_120_fu_35932_p3;
wire   [31:0] select_ln350_60_fu_35940_p3;
wire  signed [31:0] lhs_52_fu_35132_p3;
wire  signed [31:0] rhs_61_fu_32467_p3;
wire  signed [32:0] sext_ln813_114_fu_35960_p1;
wire  signed [32:0] sext_ln813_113_fu_35956_p1;
wire   [32:0] ret_V_61_fu_35964_p2;
wire   [31:0] p_Val2_363_fu_35978_p2;
wire   [0:0] p_Result_363_fu_35970_p3;
wire   [0:0] p_Result_364_fu_35984_p3;
wire   [0:0] xor_ln895_223_fu_35992_p2;
wire   [0:0] xor_ln896_223_fu_36004_p2;
wire   [0:0] xor_ln302_122_fu_36016_p2;
wire   [0:0] overflow_142_fu_35998_p2;
wire   [0:0] xor_ln302_123_fu_36022_p2;
wire   [0:0] underflow_142_fu_36010_p2;
wire   [0:0] or_ln302_61_fu_36028_p2;
wire   [31:0] select_ln302_122_fu_36034_p3;
wire   [31:0] select_ln350_61_fu_36042_p3;
wire  signed [31:0] lhs_53_fu_35234_p3;
wire  signed [31:0] rhs_62_fu_32615_p3;
wire  signed [32:0] sext_ln813_116_fu_36062_p1;
wire  signed [32:0] sext_ln813_115_fu_36058_p1;
wire   [32:0] ret_V_62_fu_36066_p2;
wire   [31:0] p_Val2_365_fu_36080_p2;
wire   [0:0] p_Result_365_fu_36072_p3;
wire   [0:0] p_Result_366_fu_36086_p3;
wire   [0:0] xor_ln895_224_fu_36094_p2;
wire   [0:0] xor_ln896_224_fu_36106_p2;
wire   [0:0] xor_ln302_124_fu_36118_p2;
wire   [0:0] overflow_143_fu_36100_p2;
wire   [0:0] xor_ln302_125_fu_36124_p2;
wire   [0:0] underflow_143_fu_36112_p2;
wire   [0:0] or_ln302_62_fu_36130_p2;
wire   [31:0] select_ln302_124_fu_36136_p3;
wire   [31:0] select_ln350_62_fu_36144_p3;
wire   [0:0] xor_ln896_126_fu_36163_p2;
wire   [0:0] xor_ln888_123_fu_36173_p2;
wire   [0:0] or_ln888_63_fu_36178_p2;
wire   [0:0] tmp_375_fu_36188_p3;
wire   [0:0] xor_ln890_61_fu_36196_p2;
wire   [0:0] or_ln890_63_fu_36202_p2;
wire   [0:0] carry_124_fu_36168_p2;
wire   [0:0] deleted_zeros_60_fu_36183_p2;
wire   [0:0] xor_ln895_126_fu_36218_p2;
wire   [0:0] or_ln895_63_fu_36224_p2;
wire   [0:0] xor_ln895_127_fu_36229_p2;
wire   [0:0] deleted_ones_63_fu_36208_p2;
wire   [0:0] xor_ln896_127_fu_36240_p2;
wire   [0:0] and_ln891_63_fu_36213_p2;
wire   [0:0] or_ln896_63_fu_36246_p2;
wire   [0:0] xor_ln896_306_fu_36252_p2;
wire   [0:0] overflow_63_fu_36234_p2;
wire   [0:0] underflow_63_fu_36258_p2;
wire   [0:0] or_ln346_63_fu_36271_p2;
wire   [31:0] select_ln346_126_fu_36263_p3;
wire  signed [31:0] sext_ln856_60_fu_36160_p1;
wire   [0:0] xor_ln896_128_fu_36288_p2;
wire   [0:0] xor_ln888_125_fu_36298_p2;
wire   [0:0] or_ln888_64_fu_36303_p2;
wire   [0:0] tmp_381_fu_36313_p3;
wire   [0:0] xor_ln890_62_fu_36321_p2;
wire   [0:0] or_ln890_64_fu_36327_p2;
wire   [0:0] carry_126_fu_36293_p2;
wire   [0:0] deleted_zeros_61_fu_36308_p2;
wire   [0:0] xor_ln895_128_fu_36343_p2;
wire   [0:0] or_ln895_64_fu_36349_p2;
wire   [0:0] xor_ln895_129_fu_36354_p2;
wire   [0:0] deleted_ones_64_fu_36333_p2;
wire   [0:0] xor_ln896_129_fu_36365_p2;
wire   [0:0] and_ln891_64_fu_36338_p2;
wire   [0:0] or_ln896_64_fu_36371_p2;
wire   [0:0] xor_ln896_307_fu_36377_p2;
wire   [0:0] overflow_64_fu_36359_p2;
wire   [0:0] underflow_64_fu_36383_p2;
wire   [0:0] or_ln346_64_fu_36396_p2;
wire   [31:0] select_ln346_128_fu_36388_p3;
wire  signed [31:0] sext_ln856_61_fu_36285_p1;
wire   [0:0] xor_ln896_130_fu_36413_p2;
wire   [0:0] xor_ln888_127_fu_36423_p2;
wire   [0:0] or_ln888_65_fu_36428_p2;
wire   [0:0] tmp_387_fu_36438_p3;
wire   [0:0] xor_ln890_63_fu_36446_p2;
wire   [0:0] or_ln890_65_fu_36452_p2;
wire   [0:0] carry_128_fu_36418_p2;
wire   [0:0] deleted_zeros_62_fu_36433_p2;
wire   [0:0] xor_ln895_130_fu_36468_p2;
wire   [0:0] or_ln895_65_fu_36474_p2;
wire   [0:0] xor_ln895_131_fu_36479_p2;
wire   [0:0] deleted_ones_65_fu_36458_p2;
wire   [0:0] xor_ln896_131_fu_36490_p2;
wire   [0:0] and_ln891_65_fu_36463_p2;
wire   [0:0] or_ln896_65_fu_36496_p2;
wire   [0:0] xor_ln896_308_fu_36502_p2;
wire   [0:0] overflow_65_fu_36484_p2;
wire   [0:0] underflow_65_fu_36508_p2;
wire   [0:0] or_ln346_65_fu_36521_p2;
wire   [31:0] select_ln346_130_fu_36513_p3;
wire  signed [31:0] sext_ln856_62_fu_36410_p1;
wire   [0:0] xor_ln896_132_fu_36538_p2;
wire   [0:0] xor_ln888_129_fu_36548_p2;
wire   [0:0] or_ln888_66_fu_36553_p2;
wire   [0:0] tmp_393_fu_36563_p3;
wire   [0:0] xor_ln890_64_fu_36571_p2;
wire   [0:0] or_ln890_66_fu_36577_p2;
wire   [0:0] carry_130_fu_36543_p2;
wire   [0:0] deleted_zeros_63_fu_36558_p2;
wire   [0:0] xor_ln895_132_fu_36593_p2;
wire   [0:0] or_ln895_66_fu_36599_p2;
wire   [0:0] xor_ln895_133_fu_36604_p2;
wire   [0:0] deleted_ones_66_fu_36583_p2;
wire   [0:0] xor_ln896_133_fu_36615_p2;
wire   [0:0] and_ln891_66_fu_36588_p2;
wire   [0:0] or_ln896_66_fu_36621_p2;
wire   [0:0] xor_ln896_309_fu_36627_p2;
wire   [0:0] overflow_66_fu_36609_p2;
wire   [0:0] underflow_66_fu_36633_p2;
wire   [0:0] or_ln346_66_fu_36646_p2;
wire   [31:0] select_ln346_132_fu_36638_p3;
wire  signed [31:0] sext_ln856_63_fu_36535_p1;
wire   [0:0] xor_ln896_134_fu_36663_p2;
wire   [0:0] xor_ln888_131_fu_36673_p2;
wire   [0:0] or_ln888_67_fu_36678_p2;
wire   [0:0] tmp_399_fu_36688_p3;
wire   [0:0] xor_ln890_65_fu_36696_p2;
wire   [0:0] or_ln890_67_fu_36702_p2;
wire   [0:0] carry_132_fu_36668_p2;
wire   [0:0] deleted_zeros_64_fu_36683_p2;
wire   [0:0] xor_ln895_134_fu_36718_p2;
wire   [0:0] or_ln895_67_fu_36724_p2;
wire   [0:0] xor_ln895_135_fu_36729_p2;
wire   [0:0] deleted_ones_67_fu_36708_p2;
wire   [0:0] xor_ln896_135_fu_36740_p2;
wire   [0:0] and_ln891_67_fu_36713_p2;
wire   [0:0] or_ln896_67_fu_36746_p2;
wire   [0:0] xor_ln896_310_fu_36752_p2;
wire   [0:0] overflow_67_fu_36734_p2;
wire   [0:0] underflow_67_fu_36758_p2;
wire   [0:0] or_ln346_67_fu_36771_p2;
wire   [31:0] select_ln346_134_fu_36763_p3;
wire  signed [31:0] sext_ln856_64_fu_36660_p1;
wire   [31:0] select_ln346_136_fu_36788_p3;
wire  signed [31:0] sext_ln856_65_fu_36785_p1;
wire   [0:0] xor_ln896_138_fu_36805_p2;
wire   [0:0] xor_ln888_135_fu_36815_p2;
wire   [0:0] or_ln888_69_fu_36820_p2;
wire   [0:0] tmp_411_fu_36830_p3;
wire   [0:0] xor_ln890_67_fu_36838_p2;
wire   [0:0] or_ln890_69_fu_36844_p2;
wire   [0:0] carry_136_fu_36810_p2;
wire   [0:0] deleted_zeros_66_fu_36825_p2;
wire   [0:0] xor_ln895_138_fu_36860_p2;
wire   [0:0] or_ln895_69_fu_36866_p2;
wire   [0:0] xor_ln895_139_fu_36871_p2;
wire   [0:0] deleted_ones_69_fu_36850_p2;
wire   [0:0] xor_ln896_139_fu_36882_p2;
wire   [0:0] and_ln891_69_fu_36855_p2;
wire   [0:0] or_ln896_69_fu_36888_p2;
wire   [0:0] xor_ln896_312_fu_36894_p2;
wire   [0:0] overflow_69_fu_36876_p2;
wire   [0:0] underflow_69_fu_36900_p2;
wire   [0:0] or_ln346_69_fu_36913_p2;
wire   [31:0] select_ln346_138_fu_36905_p3;
wire  signed [31:0] sext_ln856_66_fu_36802_p1;
wire   [0:0] xor_ln896_140_fu_36930_p2;
wire   [0:0] xor_ln888_137_fu_36940_p2;
wire   [0:0] or_ln888_70_fu_36945_p2;
wire   [0:0] tmp_417_fu_36955_p3;
wire   [0:0] xor_ln890_68_fu_36963_p2;
wire   [0:0] or_ln890_70_fu_36969_p2;
wire   [0:0] carry_138_fu_36935_p2;
wire   [0:0] deleted_zeros_67_fu_36950_p2;
wire   [0:0] xor_ln895_140_fu_36985_p2;
wire   [0:0] or_ln895_70_fu_36991_p2;
wire   [0:0] xor_ln895_141_fu_36996_p2;
wire   [0:0] deleted_ones_70_fu_36975_p2;
wire   [0:0] xor_ln896_141_fu_37007_p2;
wire   [0:0] and_ln891_70_fu_36980_p2;
wire   [0:0] or_ln896_70_fu_37013_p2;
wire   [0:0] xor_ln896_313_fu_37019_p2;
wire   [0:0] overflow_70_fu_37001_p2;
wire   [0:0] underflow_70_fu_37025_p2;
wire   [0:0] or_ln346_70_fu_37038_p2;
wire   [31:0] select_ln346_140_fu_37030_p3;
wire  signed [31:0] sext_ln856_67_fu_36927_p1;
wire   [0:0] xor_ln896_142_fu_37055_p2;
wire   [0:0] xor_ln888_139_fu_37065_p2;
wire   [0:0] or_ln888_71_fu_37070_p2;
wire   [0:0] tmp_423_fu_37080_p3;
wire   [0:0] xor_ln890_69_fu_37088_p2;
wire   [0:0] or_ln890_71_fu_37094_p2;
wire   [0:0] carry_140_fu_37060_p2;
wire   [0:0] deleted_zeros_68_fu_37075_p2;
wire   [0:0] xor_ln895_142_fu_37110_p2;
wire   [0:0] or_ln895_71_fu_37116_p2;
wire   [0:0] xor_ln895_143_fu_37121_p2;
wire   [0:0] deleted_ones_71_fu_37100_p2;
wire   [0:0] xor_ln896_143_fu_37132_p2;
wire   [0:0] and_ln891_71_fu_37105_p2;
wire   [0:0] or_ln896_71_fu_37138_p2;
wire   [0:0] xor_ln896_314_fu_37144_p2;
wire   [0:0] overflow_71_fu_37126_p2;
wire   [0:0] underflow_71_fu_37150_p2;
wire   [0:0] or_ln346_71_fu_37163_p2;
wire   [31:0] select_ln346_142_fu_37155_p3;
wire  signed [31:0] sext_ln856_68_fu_37052_p1;
wire   [20:0] zext_ln377_72_fu_37180_p1;
wire  signed [20:0] sext_ln823_69_fu_37177_p1;
wire  signed [20:0] p_Val2_215_fu_37183_p2;
wire   [0:0] p_Result_216_fu_37193_p3;
wire   [0:0] xor_ln896_144_fu_37201_p2;
wire   [0:0] xor_ln888_141_fu_37212_p2;
wire   [0:0] or_ln888_72_fu_37217_p2;
wire   [0:0] tmp_429_fu_37228_p3;
wire   [0:0] xor_ln890_70_fu_37236_p2;
wire   [0:0] or_ln890_72_fu_37242_p2;
wire   [0:0] carry_142_fu_37207_p2;
wire   [0:0] deleted_zeros_69_fu_37223_p2;
wire   [0:0] xor_ln895_144_fu_37258_p2;
wire   [0:0] or_ln895_72_fu_37264_p2;
wire   [0:0] xor_ln895_145_fu_37270_p2;
wire   [0:0] deleted_ones_72_fu_37248_p2;
wire   [0:0] xor_ln896_145_fu_37281_p2;
wire   [0:0] and_ln891_72_fu_37253_p2;
wire   [0:0] or_ln896_72_fu_37287_p2;
wire   [0:0] xor_ln896_315_fu_37293_p2;
wire   [0:0] overflow_72_fu_37275_p2;
wire   [0:0] underflow_72_fu_37299_p2;
wire   [0:0] or_ln346_72_fu_37312_p2;
wire   [31:0] select_ln346_144_fu_37304_p3;
wire  signed [31:0] sext_ln856_69_fu_37189_p1;
wire   [19:0] zext_ln377_73_fu_37329_p1;
wire  signed [19:0] sext_ln823_70_fu_37326_p1;
wire  signed [19:0] p_Val2_218_fu_37332_p2;
wire   [0:0] p_Result_219_fu_37342_p3;
wire   [0:0] xor_ln896_146_fu_37350_p2;
wire   [0:0] xor_ln888_143_fu_37361_p2;
wire   [0:0] or_ln888_73_fu_37366_p2;
wire   [0:0] tmp_435_fu_37377_p3;
wire   [0:0] xor_ln890_71_fu_37385_p2;
wire   [0:0] or_ln890_73_fu_37391_p2;
wire   [0:0] carry_144_fu_37356_p2;
wire   [0:0] deleted_zeros_70_fu_37372_p2;
wire   [0:0] xor_ln895_146_fu_37407_p2;
wire   [0:0] or_ln895_73_fu_37413_p2;
wire   [0:0] xor_ln895_147_fu_37419_p2;
wire   [0:0] deleted_ones_73_fu_37397_p2;
wire   [0:0] xor_ln896_147_fu_37430_p2;
wire   [0:0] and_ln891_73_fu_37402_p2;
wire   [0:0] or_ln896_73_fu_37436_p2;
wire   [0:0] xor_ln896_316_fu_37442_p2;
wire   [0:0] overflow_73_fu_37424_p2;
wire   [0:0] underflow_73_fu_37448_p2;
wire   [0:0] or_ln346_73_fu_37461_p2;
wire   [31:0] select_ln346_146_fu_37453_p3;
wire  signed [31:0] sext_ln856_70_fu_37338_p1;
wire   [18:0] zext_ln377_74_fu_37478_p1;
wire  signed [18:0] sext_ln823_71_fu_37475_p1;
wire  signed [18:0] p_Val2_221_fu_37481_p2;
wire   [0:0] p_Result_222_fu_37491_p3;
wire   [0:0] xor_ln896_148_fu_37499_p2;
wire   [0:0] xor_ln888_145_fu_37510_p2;
wire   [0:0] or_ln888_74_fu_37515_p2;
wire   [0:0] tmp_441_fu_37526_p3;
wire   [0:0] xor_ln890_72_fu_37534_p2;
wire   [0:0] or_ln890_74_fu_37540_p2;
wire   [0:0] carry_146_fu_37505_p2;
wire   [0:0] deleted_zeros_71_fu_37521_p2;
wire   [0:0] xor_ln895_148_fu_37556_p2;
wire   [0:0] or_ln895_74_fu_37562_p2;
wire   [0:0] xor_ln895_149_fu_37568_p2;
wire   [0:0] deleted_ones_74_fu_37546_p2;
wire   [0:0] xor_ln896_149_fu_37579_p2;
wire   [0:0] and_ln891_74_fu_37551_p2;
wire   [0:0] or_ln896_74_fu_37585_p2;
wire   [0:0] xor_ln896_317_fu_37591_p2;
wire   [0:0] overflow_74_fu_37573_p2;
wire   [0:0] underflow_74_fu_37597_p2;
wire   [0:0] or_ln346_74_fu_37610_p2;
wire   [31:0] select_ln346_148_fu_37602_p3;
wire  signed [31:0] sext_ln856_71_fu_37487_p1;
wire   [19:0] zext_ln377_75_fu_37627_p1;
wire  signed [19:0] sext_ln823_72_fu_37624_p1;
wire  signed [19:0] p_Val2_224_fu_37630_p2;
wire   [0:0] p_Result_225_fu_37640_p3;
wire   [0:0] xor_ln896_150_fu_37648_p2;
wire   [0:0] xor_ln888_147_fu_37659_p2;
wire   [0:0] or_ln888_75_fu_37664_p2;
wire   [0:0] tmp_447_fu_37675_p3;
wire   [0:0] xor_ln890_73_fu_37683_p2;
wire   [0:0] or_ln890_75_fu_37689_p2;
wire   [0:0] carry_148_fu_37654_p2;
wire   [0:0] deleted_zeros_72_fu_37670_p2;
wire   [0:0] xor_ln895_150_fu_37705_p2;
wire   [0:0] or_ln895_75_fu_37711_p2;
wire   [0:0] xor_ln895_151_fu_37717_p2;
wire   [0:0] deleted_ones_75_fu_37695_p2;
wire   [0:0] xor_ln896_151_fu_37728_p2;
wire   [0:0] and_ln891_75_fu_37700_p2;
wire   [0:0] or_ln896_75_fu_37734_p2;
wire   [0:0] xor_ln896_318_fu_37740_p2;
wire   [0:0] overflow_75_fu_37722_p2;
wire   [0:0] underflow_75_fu_37746_p2;
wire   [0:0] or_ln346_75_fu_37759_p2;
wire   [31:0] select_ln346_150_fu_37751_p3;
wire  signed [31:0] sext_ln856_72_fu_37636_p1;
wire   [31:0] select_ln346_152_fu_37776_p3;
wire  signed [31:0] sext_ln856_73_fu_37773_p1;
wire   [17:0] zext_ln377_77_fu_37793_p1;
wire  signed [17:0] sext_ln823_74_fu_37790_p1;
wire  signed [17:0] p_Val2_230_fu_37796_p2;
wire   [0:0] p_Result_231_fu_37806_p3;
wire   [0:0] xor_ln896_154_fu_37814_p2;
wire   [0:0] xor_ln888_151_fu_37825_p2;
wire   [0:0] or_ln888_77_fu_37830_p2;
wire   [0:0] tmp_459_fu_37841_p3;
wire   [0:0] xor_ln890_75_fu_37849_p2;
wire   [0:0] or_ln890_77_fu_37855_p2;
wire   [0:0] carry_152_fu_37820_p2;
wire   [0:0] deleted_zeros_74_fu_37836_p2;
wire   [0:0] xor_ln895_154_fu_37871_p2;
wire   [0:0] or_ln895_77_fu_37877_p2;
wire   [0:0] xor_ln895_155_fu_37883_p2;
wire   [0:0] deleted_ones_77_fu_37861_p2;
wire   [0:0] xor_ln896_155_fu_37894_p2;
wire   [0:0] and_ln891_77_fu_37866_p2;
wire   [0:0] or_ln896_77_fu_37900_p2;
wire   [0:0] xor_ln896_320_fu_37906_p2;
wire   [0:0] overflow_77_fu_37888_p2;
wire   [0:0] underflow_77_fu_37912_p2;
wire   [0:0] or_ln346_77_fu_37925_p2;
wire   [31:0] select_ln346_154_fu_37917_p3;
wire  signed [31:0] sext_ln856_74_fu_37802_p1;
wire   [16:0] zext_ln377_78_fu_37942_p1;
wire  signed [16:0] sext_ln823_75_fu_37939_p1;
wire  signed [16:0] p_Val2_233_fu_37945_p2;
wire   [0:0] p_Result_234_fu_37955_p3;
wire   [0:0] xor_ln896_156_fu_37963_p2;
wire   [0:0] xor_ln888_153_fu_37974_p2;
wire   [0:0] or_ln888_78_fu_37979_p2;
wire   [0:0] tmp_465_fu_37990_p3;
wire   [0:0] xor_ln890_76_fu_37998_p2;
wire   [0:0] or_ln890_78_fu_38004_p2;
wire   [0:0] carry_154_fu_37969_p2;
wire   [0:0] deleted_zeros_75_fu_37985_p2;
wire   [0:0] xor_ln895_156_fu_38020_p2;
wire   [0:0] or_ln895_78_fu_38026_p2;
wire   [0:0] xor_ln895_157_fu_38032_p2;
wire   [0:0] deleted_ones_78_fu_38010_p2;
wire   [0:0] xor_ln896_157_fu_38043_p2;
wire   [0:0] and_ln891_78_fu_38015_p2;
wire   [0:0] or_ln896_78_fu_38049_p2;
wire   [0:0] xor_ln896_321_fu_38055_p2;
wire   [0:0] overflow_78_fu_38037_p2;
wire   [0:0] underflow_78_fu_38061_p2;
wire   [0:0] or_ln346_78_fu_38074_p2;
wire   [31:0] select_ln346_156_fu_38066_p3;
wire  signed [31:0] sext_ln856_75_fu_37951_p1;
wire   [22:0] zext_ln377_79_fu_38091_p1;
wire  signed [22:0] sext_ln823_76_fu_38088_p1;
wire  signed [22:0] p_Val2_236_fu_38094_p2;
wire   [0:0] p_Result_237_fu_38104_p3;
wire   [0:0] xor_ln896_158_fu_38112_p2;
wire   [0:0] xor_ln888_155_fu_38123_p2;
wire   [0:0] or_ln888_79_fu_38128_p2;
wire   [0:0] tmp_471_fu_38139_p3;
wire   [0:0] xor_ln890_77_fu_38147_p2;
wire   [0:0] or_ln890_79_fu_38153_p2;
wire   [0:0] carry_156_fu_38118_p2;
wire   [0:0] deleted_zeros_76_fu_38134_p2;
wire   [0:0] xor_ln895_158_fu_38169_p2;
wire   [0:0] or_ln895_79_fu_38175_p2;
wire   [0:0] xor_ln895_159_fu_38181_p2;
wire   [0:0] deleted_ones_79_fu_38159_p2;
wire   [0:0] xor_ln896_159_fu_38192_p2;
wire   [0:0] and_ln891_79_fu_38164_p2;
wire   [0:0] or_ln896_79_fu_38198_p2;
wire   [0:0] xor_ln896_322_fu_38204_p2;
wire   [0:0] overflow_79_fu_38186_p2;
wire   [0:0] underflow_79_fu_38210_p2;
wire   [0:0] or_ln346_79_fu_38223_p2;
wire   [31:0] select_ln346_158_fu_38215_p3;
wire  signed [31:0] sext_ln856_76_fu_38100_p1;
wire   [30:0] zext_ln377_80_fu_38240_p1;
wire  signed [30:0] sext_ln823_77_fu_38237_p1;
wire  signed [30:0] p_Val2_239_fu_38243_p2;
wire   [0:0] p_Result_240_fu_38253_p3;
wire   [0:0] xor_ln896_160_fu_38261_p2;
wire   [0:0] xor_ln888_157_fu_38272_p2;
wire   [0:0] or_ln888_80_fu_38277_p2;
wire   [0:0] tmp_477_fu_38288_p3;
wire   [0:0] xor_ln890_78_fu_38296_p2;
wire   [0:0] or_ln890_80_fu_38302_p2;
wire   [0:0] carry_158_fu_38267_p2;
wire   [0:0] deleted_zeros_77_fu_38283_p2;
wire   [0:0] xor_ln895_160_fu_38318_p2;
wire   [0:0] or_ln895_80_fu_38324_p2;
wire   [0:0] xor_ln895_161_fu_38330_p2;
wire   [0:0] deleted_ones_80_fu_38308_p2;
wire   [0:0] xor_ln896_161_fu_38341_p2;
wire   [0:0] and_ln891_80_fu_38313_p2;
wire   [0:0] or_ln896_80_fu_38347_p2;
wire   [0:0] xor_ln896_323_fu_38353_p2;
wire   [0:0] overflow_80_fu_38335_p2;
wire   [0:0] underflow_80_fu_38359_p2;
wire   [0:0] or_ln346_80_fu_38372_p2;
wire   [31:0] select_ln346_160_fu_38364_p3;
wire  signed [31:0] sext_ln856_77_fu_38249_p1;
wire  signed [31:0] rhs_63_fu_36277_p3;
wire  signed [32:0] sext_ln813_118_fu_38389_p1;
wire  signed [32:0] sext_ln813_117_fu_38386_p1;
wire   [32:0] ret_V_63_fu_38393_p2;
wire   [31:0] p_Val2_367_fu_38407_p2;
wire   [0:0] p_Result_367_fu_38399_p3;
wire   [0:0] p_Result_368_fu_38412_p3;
wire   [0:0] xor_ln895_225_fu_38420_p2;
wire   [0:0] xor_ln896_225_fu_38432_p2;
wire   [0:0] xor_ln302_126_fu_38444_p2;
wire   [0:0] overflow_144_fu_38426_p2;
wire   [0:0] xor_ln302_127_fu_38450_p2;
wire   [0:0] underflow_144_fu_38438_p2;
wire   [0:0] or_ln302_63_fu_38456_p2;
wire   [31:0] select_ln302_126_fu_38462_p3;
wire   [31:0] select_ln350_63_fu_38470_p3;
wire  signed [31:0] rhs_64_fu_36402_p3;
wire  signed [32:0] sext_ln813_120_fu_38489_p1;
wire  signed [32:0] sext_ln813_119_fu_38486_p1;
wire   [32:0] ret_V_64_fu_38493_p2;
wire   [31:0] p_Val2_369_fu_38507_p2;
wire   [0:0] p_Result_369_fu_38499_p3;
wire   [0:0] p_Result_370_fu_38512_p3;
wire   [0:0] xor_ln895_226_fu_38520_p2;
wire   [0:0] xor_ln896_226_fu_38532_p2;
wire   [0:0] xor_ln302_128_fu_38544_p2;
wire   [0:0] overflow_145_fu_38526_p2;
wire   [0:0] xor_ln302_129_fu_38550_p2;
wire   [0:0] underflow_145_fu_38538_p2;
wire   [0:0] or_ln302_64_fu_38556_p2;
wire   [31:0] select_ln302_128_fu_38562_p3;
wire   [31:0] select_ln350_64_fu_38570_p3;
wire  signed [31:0] rhs_65_fu_36527_p3;
wire  signed [32:0] sext_ln813_122_fu_38589_p1;
wire  signed [32:0] sext_ln813_121_fu_38586_p1;
wire   [32:0] ret_V_65_fu_38593_p2;
wire   [31:0] p_Val2_371_fu_38607_p2;
wire   [0:0] p_Result_371_fu_38599_p3;
wire   [0:0] p_Result_372_fu_38612_p3;
wire   [0:0] xor_ln895_227_fu_38620_p2;
wire   [0:0] xor_ln896_227_fu_38632_p2;
wire   [0:0] xor_ln302_130_fu_38644_p2;
wire   [0:0] overflow_146_fu_38626_p2;
wire   [0:0] xor_ln302_131_fu_38650_p2;
wire   [0:0] underflow_146_fu_38638_p2;
wire   [0:0] or_ln302_65_fu_38656_p2;
wire   [31:0] select_ln302_130_fu_38662_p3;
wire   [31:0] select_ln350_65_fu_38670_p3;
wire  signed [31:0] rhs_66_fu_36652_p3;
wire  signed [32:0] sext_ln813_124_fu_38689_p1;
wire  signed [32:0] sext_ln813_123_fu_38686_p1;
wire   [32:0] ret_V_66_fu_38693_p2;
wire   [31:0] p_Val2_373_fu_38707_p2;
wire   [0:0] p_Result_373_fu_38699_p3;
wire   [0:0] p_Result_374_fu_38712_p3;
wire   [0:0] xor_ln895_228_fu_38720_p2;
wire   [0:0] xor_ln896_228_fu_38732_p2;
wire   [0:0] xor_ln302_132_fu_38744_p2;
wire   [0:0] overflow_147_fu_38726_p2;
wire   [0:0] xor_ln302_133_fu_38750_p2;
wire   [0:0] underflow_147_fu_38738_p2;
wire   [0:0] or_ln302_66_fu_38756_p2;
wire   [31:0] select_ln302_132_fu_38762_p3;
wire   [31:0] select_ln350_66_fu_38770_p3;
wire  signed [31:0] rhs_67_fu_36777_p3;
wire  signed [32:0] sext_ln813_126_fu_38789_p1;
wire  signed [32:0] sext_ln813_125_fu_38786_p1;
wire   [32:0] ret_V_67_fu_38793_p2;
wire   [31:0] p_Val2_375_fu_38807_p2;
wire   [0:0] p_Result_375_fu_38799_p3;
wire   [0:0] p_Result_376_fu_38812_p3;
wire   [0:0] xor_ln895_229_fu_38820_p2;
wire   [0:0] xor_ln896_229_fu_38832_p2;
wire   [0:0] xor_ln302_134_fu_38844_p2;
wire   [0:0] overflow_148_fu_38826_p2;
wire   [0:0] xor_ln302_135_fu_38850_p2;
wire   [0:0] underflow_148_fu_38838_p2;
wire   [0:0] or_ln302_67_fu_38856_p2;
wire   [31:0] select_ln302_134_fu_38862_p3;
wire   [31:0] select_ln350_67_fu_38870_p3;
wire  signed [31:0] rhs_68_fu_36795_p3;
wire  signed [32:0] sext_ln813_128_fu_38889_p1;
wire  signed [32:0] sext_ln813_127_fu_38886_p1;
wire   [32:0] ret_V_68_fu_38893_p2;
wire   [31:0] p_Val2_377_fu_38907_p2;
wire   [0:0] p_Result_377_fu_38899_p3;
wire   [0:0] p_Result_378_fu_38912_p3;
wire   [0:0] xor_ln895_230_fu_38920_p2;
wire   [0:0] xor_ln896_230_fu_38932_p2;
wire   [0:0] xor_ln302_136_fu_38944_p2;
wire   [0:0] overflow_149_fu_38926_p2;
wire   [0:0] xor_ln302_137_fu_38950_p2;
wire   [0:0] underflow_149_fu_38938_p2;
wire   [0:0] or_ln302_68_fu_38956_p2;
wire   [31:0] select_ln302_136_fu_38962_p3;
wire   [31:0] select_ln350_68_fu_38970_p3;
wire  signed [31:0] rhs_69_fu_36919_p3;
wire  signed [32:0] sext_ln813_130_fu_38989_p1;
wire  signed [32:0] sext_ln813_129_fu_38986_p1;
wire   [32:0] ret_V_69_fu_38993_p2;
wire   [31:0] p_Val2_379_fu_39007_p2;
wire   [0:0] p_Result_379_fu_38999_p3;
wire   [0:0] p_Result_380_fu_39012_p3;
wire   [0:0] xor_ln895_231_fu_39020_p2;
wire   [0:0] xor_ln896_231_fu_39032_p2;
wire   [0:0] xor_ln302_138_fu_39044_p2;
wire   [0:0] overflow_150_fu_39026_p2;
wire   [0:0] xor_ln302_139_fu_39050_p2;
wire   [0:0] underflow_150_fu_39038_p2;
wire   [0:0] or_ln302_69_fu_39056_p2;
wire   [31:0] select_ln302_138_fu_39062_p3;
wire   [31:0] select_ln350_69_fu_39070_p3;
wire  signed [31:0] rhs_70_fu_37044_p3;
wire  signed [32:0] sext_ln813_132_fu_39089_p1;
wire  signed [32:0] sext_ln813_131_fu_39086_p1;
wire   [32:0] ret_V_70_fu_39093_p2;
wire   [31:0] p_Val2_381_fu_39107_p2;
wire   [0:0] p_Result_381_fu_39099_p3;
wire   [0:0] p_Result_382_fu_39112_p3;
wire   [0:0] xor_ln895_232_fu_39120_p2;
wire   [0:0] xor_ln896_232_fu_39132_p2;
wire   [0:0] xor_ln302_140_fu_39144_p2;
wire   [0:0] overflow_151_fu_39126_p2;
wire   [0:0] xor_ln302_141_fu_39150_p2;
wire   [0:0] underflow_151_fu_39138_p2;
wire   [0:0] or_ln302_70_fu_39156_p2;
wire   [31:0] select_ln302_140_fu_39162_p3;
wire   [31:0] select_ln350_70_fu_39170_p3;
wire  signed [31:0] rhs_71_fu_37169_p3;
wire  signed [32:0] sext_ln813_134_fu_39189_p1;
wire  signed [32:0] sext_ln813_133_fu_39186_p1;
wire   [32:0] ret_V_71_fu_39193_p2;
wire   [31:0] p_Val2_383_fu_39207_p2;
wire   [0:0] p_Result_383_fu_39199_p3;
wire   [0:0] p_Result_384_fu_39212_p3;
wire   [0:0] xor_ln895_233_fu_39220_p2;
wire   [0:0] xor_ln896_233_fu_39232_p2;
wire   [0:0] xor_ln302_142_fu_39244_p2;
wire   [0:0] overflow_152_fu_39226_p2;
wire   [0:0] xor_ln302_143_fu_39250_p2;
wire   [0:0] underflow_152_fu_39238_p2;
wire   [0:0] or_ln302_71_fu_39256_p2;
wire   [31:0] select_ln302_142_fu_39262_p3;
wire   [31:0] select_ln350_71_fu_39270_p3;
wire  signed [31:0] lhs_63_fu_38478_p3;
wire  signed [31:0] rhs_72_fu_37318_p3;
wire  signed [32:0] sext_ln813_136_fu_39290_p1;
wire  signed [32:0] sext_ln813_135_fu_39286_p1;
wire   [32:0] ret_V_72_fu_39294_p2;
wire   [31:0] p_Val2_385_fu_39308_p2;
wire   [0:0] p_Result_385_fu_39300_p3;
wire   [0:0] p_Result_386_fu_39314_p3;
wire   [0:0] xor_ln895_234_fu_39322_p2;
wire   [0:0] xor_ln896_234_fu_39334_p2;
wire   [0:0] xor_ln302_144_fu_39346_p2;
wire   [0:0] overflow_153_fu_39328_p2;
wire   [0:0] xor_ln302_145_fu_39352_p2;
wire   [0:0] underflow_153_fu_39340_p2;
wire   [0:0] or_ln302_72_fu_39358_p2;
wire   [31:0] select_ln302_144_fu_39364_p3;
wire   [31:0] select_ln350_72_fu_39372_p3;
wire  signed [31:0] lhs_64_fu_38578_p3;
wire  signed [31:0] rhs_73_fu_37467_p3;
wire  signed [32:0] sext_ln813_138_fu_39392_p1;
wire  signed [32:0] sext_ln813_137_fu_39388_p1;
wire   [32:0] ret_V_73_fu_39396_p2;
wire   [31:0] p_Val2_387_fu_39410_p2;
wire   [0:0] p_Result_387_fu_39402_p3;
wire   [0:0] p_Result_388_fu_39416_p3;
wire   [0:0] xor_ln895_235_fu_39424_p2;
wire   [0:0] xor_ln896_235_fu_39436_p2;
wire   [0:0] xor_ln302_146_fu_39448_p2;
wire   [0:0] overflow_154_fu_39430_p2;
wire   [0:0] xor_ln302_147_fu_39454_p2;
wire   [0:0] underflow_154_fu_39442_p2;
wire   [0:0] or_ln302_73_fu_39460_p2;
wire   [31:0] select_ln302_146_fu_39466_p3;
wire   [31:0] select_ln350_73_fu_39474_p3;
wire  signed [31:0] lhs_65_fu_38678_p3;
wire  signed [31:0] rhs_74_fu_37616_p3;
wire  signed [32:0] sext_ln813_140_fu_39494_p1;
wire  signed [32:0] sext_ln813_139_fu_39490_p1;
wire   [32:0] ret_V_74_fu_39498_p2;
wire   [31:0] p_Val2_389_fu_39512_p2;
wire   [0:0] p_Result_389_fu_39504_p3;
wire   [0:0] p_Result_390_fu_39518_p3;
wire   [0:0] xor_ln895_236_fu_39526_p2;
wire   [0:0] xor_ln896_236_fu_39538_p2;
wire   [0:0] xor_ln302_148_fu_39550_p2;
wire   [0:0] overflow_155_fu_39532_p2;
wire   [0:0] xor_ln302_149_fu_39556_p2;
wire   [0:0] underflow_155_fu_39544_p2;
wire   [0:0] or_ln302_74_fu_39562_p2;
wire   [31:0] select_ln302_148_fu_39568_p3;
wire   [31:0] select_ln350_74_fu_39576_p3;
wire  signed [31:0] lhs_66_fu_38778_p3;
wire  signed [31:0] rhs_75_fu_37765_p3;
wire  signed [32:0] sext_ln813_142_fu_39596_p1;
wire  signed [32:0] sext_ln813_141_fu_39592_p1;
wire   [32:0] ret_V_75_fu_39600_p2;
wire   [31:0] p_Val2_391_fu_39614_p2;
wire   [0:0] p_Result_391_fu_39606_p3;
wire   [0:0] p_Result_392_fu_39620_p3;
wire   [0:0] xor_ln895_237_fu_39628_p2;
wire   [0:0] xor_ln896_237_fu_39640_p2;
wire   [0:0] xor_ln302_150_fu_39652_p2;
wire   [0:0] overflow_156_fu_39634_p2;
wire   [0:0] xor_ln302_151_fu_39658_p2;
wire   [0:0] underflow_156_fu_39646_p2;
wire   [0:0] or_ln302_75_fu_39664_p2;
wire   [31:0] select_ln302_150_fu_39670_p3;
wire   [31:0] select_ln350_75_fu_39678_p3;
wire  signed [31:0] lhs_67_fu_38878_p3;
wire  signed [31:0] rhs_76_fu_37783_p3;
wire  signed [32:0] sext_ln813_144_fu_39698_p1;
wire  signed [32:0] sext_ln813_143_fu_39694_p1;
wire   [32:0] ret_V_76_fu_39702_p2;
wire   [31:0] p_Val2_393_fu_39716_p2;
wire   [0:0] p_Result_393_fu_39708_p3;
wire   [0:0] p_Result_394_fu_39722_p3;
wire   [0:0] xor_ln895_238_fu_39730_p2;
wire   [0:0] xor_ln896_238_fu_39742_p2;
wire   [0:0] xor_ln302_152_fu_39754_p2;
wire   [0:0] overflow_157_fu_39736_p2;
wire   [0:0] xor_ln302_153_fu_39760_p2;
wire   [0:0] underflow_157_fu_39748_p2;
wire   [0:0] or_ln302_76_fu_39766_p2;
wire   [31:0] select_ln302_152_fu_39772_p3;
wire   [31:0] select_ln350_76_fu_39780_p3;
wire  signed [31:0] lhs_68_fu_38978_p3;
wire  signed [31:0] rhs_77_fu_37931_p3;
wire  signed [32:0] sext_ln813_146_fu_39800_p1;
wire  signed [32:0] sext_ln813_145_fu_39796_p1;
wire   [32:0] ret_V_77_fu_39804_p2;
wire   [31:0] p_Val2_395_fu_39818_p2;
wire   [0:0] p_Result_395_fu_39810_p3;
wire   [0:0] p_Result_396_fu_39824_p3;
wire   [0:0] xor_ln895_239_fu_39832_p2;
wire   [0:0] xor_ln896_239_fu_39844_p2;
wire   [0:0] xor_ln302_154_fu_39856_p2;
wire   [0:0] overflow_158_fu_39838_p2;
wire   [0:0] xor_ln302_155_fu_39862_p2;
wire   [0:0] underflow_158_fu_39850_p2;
wire   [0:0] or_ln302_77_fu_39868_p2;
wire   [31:0] select_ln302_154_fu_39874_p3;
wire   [31:0] select_ln350_77_fu_39882_p3;
wire  signed [31:0] lhs_69_fu_39078_p3;
wire  signed [31:0] rhs_78_fu_38080_p3;
wire  signed [32:0] sext_ln813_148_fu_39902_p1;
wire  signed [32:0] sext_ln813_147_fu_39898_p1;
wire   [32:0] ret_V_78_fu_39906_p2;
wire   [31:0] p_Val2_397_fu_39920_p2;
wire   [0:0] p_Result_397_fu_39912_p3;
wire   [0:0] p_Result_398_fu_39926_p3;
wire   [0:0] xor_ln895_240_fu_39934_p2;
wire   [0:0] xor_ln896_240_fu_39946_p2;
wire   [0:0] xor_ln302_156_fu_39958_p2;
wire   [0:0] overflow_159_fu_39940_p2;
wire   [0:0] xor_ln302_157_fu_39964_p2;
wire   [0:0] underflow_159_fu_39952_p2;
wire   [0:0] or_ln302_78_fu_39970_p2;
wire   [31:0] select_ln302_156_fu_39976_p3;
wire   [31:0] select_ln350_78_fu_39984_p3;
wire  signed [31:0] lhs_70_fu_39178_p3;
wire  signed [31:0] rhs_79_fu_38229_p3;
wire  signed [32:0] sext_ln813_150_fu_40004_p1;
wire  signed [32:0] sext_ln813_149_fu_40000_p1;
wire   [32:0] ret_V_79_fu_40008_p2;
wire   [31:0] p_Val2_399_fu_40022_p2;
wire   [0:0] p_Result_399_fu_40014_p3;
wire   [0:0] p_Result_400_fu_40028_p3;
wire   [0:0] xor_ln895_241_fu_40036_p2;
wire   [0:0] xor_ln896_241_fu_40048_p2;
wire   [0:0] xor_ln302_158_fu_40060_p2;
wire   [0:0] overflow_160_fu_40042_p2;
wire   [0:0] xor_ln302_159_fu_40066_p2;
wire   [0:0] underflow_160_fu_40054_p2;
wire   [0:0] or_ln302_79_fu_40072_p2;
wire   [31:0] select_ln302_158_fu_40078_p3;
wire   [31:0] select_ln350_79_fu_40086_p3;
wire  signed [31:0] lhs_71_fu_39278_p3;
wire  signed [31:0] rhs_80_fu_38378_p3;
wire  signed [32:0] sext_ln813_152_fu_40106_p1;
wire  signed [32:0] sext_ln813_151_fu_40102_p1;
wire   [32:0] ret_V_80_fu_40110_p2;
wire   [31:0] p_Val2_401_fu_40124_p2;
wire   [0:0] p_Result_401_fu_40116_p3;
wire   [0:0] p_Result_402_fu_40130_p3;
wire   [0:0] xor_ln895_242_fu_40138_p2;
wire   [0:0] xor_ln896_242_fu_40150_p2;
wire   [0:0] xor_ln302_160_fu_40162_p2;
wire   [0:0] overflow_161_fu_40144_p2;
wire   [0:0] xor_ln302_161_fu_40168_p2;
wire   [0:0] underflow_161_fu_40156_p2;
wire   [0:0] or_ln302_80_fu_40174_p2;
wire   [31:0] select_ln302_160_fu_40180_p3;
wire   [31:0] select_ln350_80_fu_40188_p3;
wire   [31:0] select_ln302_145_fu_39380_p3;
wire   [31:0] select_ln302_147_fu_39482_p3;
wire   [31:0] select_ln302_149_fu_39584_p3;
wire   [31:0] select_ln302_151_fu_39686_p3;
wire   [31:0] select_ln302_153_fu_39788_p3;
wire   [31:0] select_ln302_155_fu_39890_p3;
wire   [31:0] select_ln302_157_fu_39992_p3;
wire   [31:0] select_ln302_159_fu_40094_p3;
wire   [31:0] select_ln302_161_fu_40196_p3;
reg    ap_ce_reg;
reg  signed [31:0] p_read_int_reg;
reg  signed [31:0] p_read1_int_reg;
reg  signed [31:0] p_read2_int_reg;
reg   [31:0] p_read3_int_reg;
reg   [31:0] p_read4_int_reg;
reg   [31:0] p_read5_int_reg;
reg   [31:0] p_read6_int_reg;
reg   [31:0] p_read7_int_reg;
reg   [31:0] p_read8_int_reg;
reg   [31:0] ap_return_0_int_reg;
reg   [31:0] ap_return_1_int_reg;
reg   [31:0] ap_return_2_int_reg;
reg   [31:0] ap_return_3_int_reg;
reg   [31:0] ap_return_4_int_reg;
reg   [31:0] ap_return_5_int_reg;
reg   [31:0] ap_return_6_int_reg;
reg   [31:0] ap_return_7_int_reg;
reg   [31:0] ap_return_8_int_reg;

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U156(
    .din0(p_read_int_reg),
    .din1(r_V_1_fu_470_p1),
    .dout(r_V_1_fu_470_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U157(
    .din0(r_V_47_fu_471_p0),
    .din1(r_V_47_fu_471_p1),
    .dout(r_V_47_fu_471_p2)
);

motorB_mul_32s_22ns_53_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 22 ),
    .dout_WIDTH( 53 ))
mul_32s_22ns_53_1_0_U158(
    .din0(p_read_22_reg_40302),
    .din1(r_V_41_fu_472_p1),
    .dout(r_V_41_fu_472_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U159(
    .din0(r_V_19_fu_473_p0),
    .din1(r_V_19_fu_473_p1),
    .dout(r_V_19_fu_473_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U160(
    .din0(r_V_60_fu_474_p0),
    .din1(r_V_60_fu_474_p1),
    .dout(r_V_60_fu_474_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U161(
    .din0(p_read_22_reg_40302),
    .din1(r_V_35_fu_476_p1),
    .dout(r_V_35_fu_476_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U162(
    .din0(r_V_62_fu_477_p0),
    .din1(r_V_62_fu_477_p1),
    .dout(r_V_62_fu_477_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U163(
    .din0(r_V_11_fu_478_p0),
    .din1(r_V_11_fu_478_p1),
    .dout(r_V_11_fu_478_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U164(
    .din0(r_V_49_fu_480_p0),
    .din1(r_V_49_fu_480_p1),
    .dout(r_V_49_fu_480_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U165(
    .din0(r_V_18_fu_481_p0),
    .din1(r_V_18_fu_481_p1),
    .dout(r_V_18_fu_481_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U166(
    .din0(r_V_15_fu_482_p0),
    .din1(r_V_15_fu_482_p1),
    .dout(r_V_15_fu_482_p2)
);

motorB_mul_32s_14ns_46_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 46 ))
mul_32s_14ns_46_1_0_U167(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_76_fu_484_p1),
    .dout(r_V_76_fu_484_p2)
);

motorB_mul_32s_10ns_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10ns_42_1_0_U168(
    .din0(p_read2_int_reg),
    .din1(r_V_17_fu_485_p1),
    .dout(r_V_17_fu_485_p2)
);

motorB_mul_32s_23ns_54_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 23 ),
    .dout_WIDTH( 54 ))
mul_32s_23ns_54_1_0_U169(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_77_fu_486_p1),
    .dout(r_V_77_fu_486_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U170(
    .din0(r_V_30_fu_488_p0),
    .din1(r_V_30_fu_488_p1),
    .dout(r_V_30_fu_488_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U171(
    .din0(p_read1_int_reg),
    .din1(r_V_12_fu_489_p1),
    .dout(r_V_12_fu_489_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U172(
    .din0(r_V_26_fu_490_p0),
    .din1(r_V_26_fu_490_p1),
    .dout(r_V_26_fu_490_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U173(
    .din0(p_read_20_reg_40279_pp0_iter1_reg),
    .din1(r_V_51_fu_491_p1),
    .dout(r_V_51_fu_491_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U174(
    .din0(p_read2_int_reg),
    .din1(r_V_16_fu_492_p1),
    .dout(r_V_16_fu_492_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U175(
    .din0(r_V_54_fu_493_p0),
    .din1(r_V_54_fu_493_p1),
    .dout(r_V_54_fu_493_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U176(
    .din0(r_V_37_fu_494_p0),
    .din1(r_V_37_fu_494_p1),
    .dout(r_V_37_fu_494_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U177(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_74_fu_495_p1),
    .dout(r_V_74_fu_495_p2)
);

motorB_mul_32s_14s_46_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 46 ))
mul_32s_14s_46_1_0_U178(
    .din0(p_read_23_reg_40314),
    .din1(r_V_31_fu_496_p1),
    .dout(r_V_31_fu_496_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U179(
    .din0(r_V_25_fu_497_p0),
    .din1(r_V_25_fu_497_p1),
    .dout(r_V_25_fu_497_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U180(
    .din0(r_V_38_fu_498_p0),
    .din1(r_V_38_fu_498_p1),
    .dout(r_V_38_fu_498_p2)
);

motorB_mul_32s_25s_56_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 25 ),
    .dout_WIDTH( 56 ))
mul_32s_25s_56_1_0_U181(
    .din0(r_V_32_fu_499_p0),
    .din1(r_V_32_fu_499_p1),
    .dout(r_V_32_fu_499_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U182(
    .din0(r_V_5_fu_500_p0),
    .din1(r_V_5_fu_500_p1),
    .dout(r_V_5_fu_500_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U183(
    .din0(r_V_13_fu_501_p0),
    .din1(r_V_13_fu_501_p1),
    .dout(r_V_13_fu_501_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U184(
    .din0(r_V_9_fu_503_p0),
    .din1(r_V_9_fu_503_p1),
    .dout(r_V_9_fu_503_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U185(
    .din0(r_V_57_fu_504_p0),
    .din1(r_V_57_fu_504_p1),
    .dout(r_V_57_fu_504_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U186(
    .din0(r_V_39_fu_505_p0),
    .din1(r_V_39_fu_505_p1),
    .dout(r_V_39_fu_505_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U187(
    .din0(p_read_21_reg_40289_pp0_iter1_reg),
    .din1(r_V_45_fu_506_p1),
    .dout(r_V_45_fu_506_p2)
);

motorB_mul_32s_25ns_56_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 25 ),
    .dout_WIDTH( 56 ))
mul_32s_25ns_56_1_0_U188(
    .din0(r_V_24_fu_508_p0),
    .din1(r_V_24_fu_508_p1),
    .dout(r_V_24_fu_508_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U189(
    .din0(r_V_34_fu_509_p0),
    .din1(r_V_34_fu_509_p1),
    .dout(r_V_34_fu_509_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U190(
    .din0(r_V_3_fu_510_p0),
    .din1(r_V_3_fu_510_p1),
    .dout(r_V_3_fu_510_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U191(
    .din0(r_V_66_fu_511_p0),
    .din1(r_V_66_fu_511_p1),
    .dout(r_V_66_fu_511_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U192(
    .din0(p_read_22_reg_40302),
    .din1(r_V_40_fu_512_p1),
    .dout(r_V_40_fu_512_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U193(
    .din0(r_V_8_fu_514_p0),
    .din1(r_V_8_fu_514_p1),
    .dout(r_V_8_fu_514_p2)
);

motorB_mul_32s_6s_38_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 38 ))
mul_32s_6s_38_1_0_U194(
    .din0(p_read2_int_reg),
    .din1(r_V_20_fu_515_p1),
    .dout(r_V_20_fu_515_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U195(
    .din0(r_V_70_fu_516_p0),
    .din1(r_V_70_fu_516_p1),
    .dout(r_V_70_fu_516_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U196(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_71_fu_517_p1),
    .dout(r_V_71_fu_517_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U197(
    .din0(r_V_23_fu_518_p0),
    .din1(r_V_23_fu_518_p1),
    .dout(r_V_23_fu_518_p2)
);

motorB_mul_32s_15s_47_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 47 ))
mul_32s_15s_47_1_0_U198(
    .din0(p_read_int_reg),
    .din1(r_V_fu_519_p1),
    .dout(r_V_fu_519_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U199(
    .din0(p_read_21_reg_40289_pp0_iter1_reg),
    .din1(r_V_44_fu_520_p1),
    .dout(r_V_44_fu_520_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U200(
    .din0(r_V_28_fu_521_p0),
    .din1(r_V_28_fu_521_p1),
    .dout(r_V_28_fu_521_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U201(
    .din0(r_V_67_fu_522_p0),
    .din1(r_V_67_fu_522_p1),
    .dout(r_V_67_fu_522_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U202(
    .din0(p_read_20_reg_40279_pp0_iter1_reg),
    .din1(r_V_52_fu_523_p1),
    .dout(r_V_52_fu_523_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U203(
    .din0(r_V_72_fu_525_p0),
    .din1(r_V_72_fu_525_p1),
    .dout(r_V_72_fu_525_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U204(
    .din0(r_V_4_fu_526_p0),
    .din1(r_V_4_fu_526_p1),
    .dout(r_V_4_fu_526_p2)
);

motorB_mul_32s_20s_51_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 20 ),
    .dout_WIDTH( 51 ))
mul_32s_20s_51_1_0_U205(
    .din0(p_read_22_reg_40302),
    .din1(r_V_33_fu_527_p1),
    .dout(r_V_33_fu_527_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U206(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_69_fu_529_p1),
    .dout(r_V_69_fu_529_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U207(
    .din0(p_read_21_reg_40289_pp0_iter1_reg),
    .din1(r_V_46_fu_530_p1),
    .dout(r_V_46_fu_530_p2)
);

motorB_mul_32s_11s_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11s_43_1_0_U208(
    .din0(r_V_43_fu_531_p0),
    .din1(r_V_43_fu_531_p1),
    .dout(r_V_43_fu_531_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U209(
    .din0(r_V_59_fu_532_p0),
    .din1(r_V_59_fu_532_p1),
    .dout(r_V_59_fu_532_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U210(
    .din0(r_V_64_fu_533_p0),
    .din1(r_V_64_fu_533_p1),
    .dout(r_V_64_fu_533_p2)
);

motorB_mul_32s_12ns_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12ns_44_1_0_U211(
    .din0(r_V_53_fu_534_p0),
    .din1(r_V_53_fu_534_p1),
    .dout(r_V_53_fu_534_p2)
);

motorB_mul_32s_13s_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13s_45_1_0_U212(
    .din0(p_read2_int_reg),
    .din1(r_V_22_fu_535_p1),
    .dout(r_V_22_fu_535_p2)
);

motorB_mul_32s_26s_57_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 26 ),
    .dout_WIDTH( 57 ))
mul_32s_26s_57_1_0_U213(
    .din0(p_read_int_reg),
    .din1(r_V_7_fu_537_p1),
    .dout(r_V_7_fu_537_p2)
);

motorB_mul_32s_9s_41_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 41 ))
mul_32s_9s_41_1_0_U214(
    .din0(r_V_29_fu_538_p0),
    .din1(r_V_29_fu_538_p1),
    .dout(r_V_29_fu_538_p2)
);

motorB_mul_32s_8ns_40_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 40 ))
mul_32s_8ns_40_1_0_U215(
    .din0(p_read_18_reg_40258_pp0_iter2_reg),
    .din1(r_V_75_fu_539_p1),
    .dout(r_V_75_fu_539_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U216(
    .din0(r_V_55_fu_540_p0),
    .din1(r_V_55_fu_540_p1),
    .dout(r_V_55_fu_540_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U217(
    .din0(r_V_27_fu_541_p0),
    .din1(r_V_27_fu_541_p1),
    .dout(r_V_27_fu_541_p2)
);

motorB_mul_32s_11ns_43_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 43 ))
mul_32s_11ns_43_1_0_U218(
    .din0(r_V_61_fu_543_p0),
    .din1(r_V_61_fu_543_p1),
    .dout(r_V_61_fu_543_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U219(
    .din0(r_V_68_fu_544_p0),
    .din1(r_V_68_fu_544_p1),
    .dout(r_V_68_fu_544_p2)
);

motorB_mul_32s_10s_42_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 42 ))
mul_32s_10s_42_1_0_U220(
    .din0(r_V_63_fu_545_p0),
    .din1(r_V_63_fu_545_p1),
    .dout(r_V_63_fu_545_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U221(
    .din0(r_V_14_fu_546_p0),
    .din1(r_V_14_fu_546_p1),
    .dout(r_V_14_fu_546_p2)
);

motorB_mul_32s_13ns_45_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 45 ))
mul_32s_13ns_45_1_0_U222(
    .din0(r_V_10_fu_548_p0),
    .din1(r_V_10_fu_548_p1),
    .dout(r_V_10_fu_548_p2)
);

motorB_mul_32s_12s_44_1_0 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 44 ))
mul_32s_12s_44_1_0_U223(
    .din0(r_V_56_fu_549_p0),
    .din1(r_V_56_fu_549_p1),
    .dout(r_V_56_fu_549_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        Range2_all_ones_11_reg_40651 <= r_V_10_fu_548_p2[32'd44];
        Range2_all_ones_12_reg_40680 <= r_V_11_fu_478_p2[32'd44];
        Range2_all_ones_13_reg_40726 <= r_V_12_fu_489_p2[32'd41];
        Range2_all_ones_14_reg_40755 <= r_V_13_fu_501_p2[32'd42];
        Range2_all_ones_15_reg_40784 <= r_V_14_fu_546_p2[32'd44];
        Range2_all_ones_16_reg_40813 <= r_V_15_fu_482_p2[32'd42];
        Range2_all_ones_17_reg_40842 <= r_V_16_fu_492_p2[32'd43];
        Range2_all_ones_18_reg_40871 <= r_V_17_fu_485_p2[32'd41];
        Range2_all_ones_19_reg_40900 <= r_V_18_fu_481_p2[32'd42];
        Range2_all_ones_1_reg_40378 <= r_V_1_fu_470_p2[32'd41];
        Range2_all_ones_20_reg_40929 <= r_V_19_fu_473_p2[32'd42];
        Range2_all_ones_21_reg_40958 <= r_V_20_fu_515_p2[32'd37];
        Range2_all_ones_23_reg_41002 <= r_V_22_fu_535_p2[32'd44];
        Range2_all_ones_24_reg_41031 <= r_V_23_fu_518_p2[32'd42];
        Range2_all_ones_25_reg_41172 <= r_V_24_fu_508_p2[32'd55];
        Range2_all_ones_26_reg_41203 <= r_V_25_fu_497_p2[32'd43];
        Range2_all_ones_27_reg_41234 <= r_V_26_fu_490_p2[32'd42];
        Range2_all_ones_28_reg_41265 <= r_V_27_fu_541_p2[32'd43];
        Range2_all_ones_29_reg_41296 <= r_V_28_fu_521_p2[32'd42];
        Range2_all_ones_30_reg_41327 <= r_V_29_fu_538_p2[32'd40];
        Range2_all_ones_31_reg_41358 <= r_V_30_fu_488_p2[32'd40];
        Range2_all_ones_32_reg_41389 <= r_V_31_fu_496_p2[32'd45];
        Range2_all_ones_33_reg_41420 <= r_V_32_fu_499_p2[32'd55];
        Range2_all_ones_34_reg_41449 <= r_V_33_fu_527_p2[32'd50];
        Range2_all_ones_35_reg_41478 <= r_V_34_fu_509_p2[32'd43];
        Range2_all_ones_36_reg_41507 <= r_V_35_fu_476_p2[32'd41];
        Range2_all_ones_38_reg_41551 <= r_V_37_fu_494_p2[32'd42];
        Range2_all_ones_39_reg_41580 <= r_V_38_fu_498_p2[32'd43];
        Range2_all_ones_3_reg_40424 <= r_V_3_fu_510_p2[32'd44];
        Range2_all_ones_40_reg_41609 <= r_V_39_fu_505_p2[32'd42];
        Range2_all_ones_41_reg_41638 <= r_V_40_fu_512_p2[32'd44];
        Range2_all_ones_42_reg_41667 <= r_V_41_fu_472_p2[32'd52];
        Range2_all_ones_44_reg_41795 <= r_V_43_fu_531_p2[32'd42];
        Range2_all_ones_45_reg_41826 <= r_V_44_fu_520_p2[32'd41];
        Range2_all_ones_46_reg_41857 <= r_V_45_fu_506_p2[32'd44];
        Range2_all_ones_47_reg_41888 <= r_V_46_fu_530_p2[32'd43];
        Range2_all_ones_48_reg_41919 <= r_V_47_fu_471_p2[32'd42];
        Range2_all_ones_4_reg_40455 <= r_V_4_fu_526_p2[32'd42];
        Range2_all_ones_50_reg_41965 <= r_V_49_fu_480_p2[32'd42];
        Range2_all_ones_52_reg_42009 <= r_V_51_fu_491_p2[32'd42];
        Range2_all_ones_53_reg_42038 <= r_V_52_fu_523_p2[32'd41];
        Range2_all_ones_54_reg_42067 <= r_V_53_fu_534_p2[32'd43];
        Range2_all_ones_55_reg_42096 <= r_V_54_fu_493_p2[32'd44];
        Range2_all_ones_56_reg_42125 <= r_V_55_fu_540_p2[32'd44];
        Range2_all_ones_57_reg_42154 <= r_V_56_fu_549_p2[32'd43];
        Range2_all_ones_58_reg_42183 <= r_V_57_fu_504_p2[32'd44];
        Range2_all_ones_5_reg_40486 <= r_V_5_fu_500_p2[32'd42];
        Range2_all_ones_60_reg_42227 <= r_V_59_fu_532_p2[32'd43];
        Range2_all_ones_61_reg_42410 <= r_V_60_fu_474_p2[32'd41];
        Range2_all_ones_62_reg_42441 <= r_V_61_fu_543_p2[32'd42];
        Range2_all_ones_63_reg_42472 <= r_V_62_fu_477_p2[32'd43];
        Range2_all_ones_64_reg_42503 <= r_V_63_fu_545_p2[32'd41];
        Range2_all_ones_65_reg_42534 <= r_V_64_fu_533_p2[32'd43];
        Range2_all_ones_67_reg_42580 <= r_V_66_fu_511_p2[32'd42];
        Range2_all_ones_68_reg_42611 <= r_V_67_fu_522_p2[32'd43];
        Range2_all_ones_69_reg_42642 <= r_V_68_fu_544_p2[32'd41];
        Range2_all_ones_70_reg_42671 <= r_V_69_fu_529_p2[32'd43];
        Range2_all_ones_71_reg_42700 <= r_V_70_fu_516_p2[32'd42];
        Range2_all_ones_72_reg_42729 <= r_V_71_fu_517_p2[32'd41];
        Range2_all_ones_73_reg_42758 <= r_V_72_fu_525_p2[32'd42];
        Range2_all_ones_75_reg_42802 <= r_V_74_fu_495_p2[32'd40];
        Range2_all_ones_76_reg_42831 <= r_V_75_fu_539_p2[32'd39];
        Range2_all_ones_77_reg_42860 <= r_V_76_fu_484_p2[32'd45];
        Range2_all_ones_78_reg_42889 <= r_V_77_fu_486_p2[32'd53];
        Range2_all_ones_7_reg_40532 <= r_V_7_fu_537_p2[32'd56];
        Range2_all_ones_8_reg_40563 <= r_V_8_fu_514_p2[32'd44];
        Range2_all_ones_9_reg_40592 <= r_V_9_fu_503_p2[32'd42];
        Range2_all_ones_reg_40347 <= r_V_fu_519_p2[32'd46];
        lhs_10_reg_41680 <= lhs_10_fu_23616_p3;
        lhs_12_reg_41686 <= lhs_12_fu_23820_p3;
        lhs_13_reg_41692 <= lhs_13_fu_23922_p3;
        lhs_14_reg_41698 <= lhs_14_fu_24024_p3;
        lhs_16_reg_41704 <= lhs_16_fu_24228_p3;
        lhs_17_reg_41710 <= lhs_17_fu_24330_p3;
        lhs_38_reg_42274 <= lhs_38_fu_30323_p3;
        lhs_42_reg_42340 <= lhs_42_fu_30533_p3;
        lhs_54_reg_42896 <= lhs_54_fu_35336_p3;
        lhs_55_reg_42902 <= lhs_55_fu_35438_p3;
        lhs_56_reg_42908 <= lhs_56_fu_35540_p3;
        lhs_57_reg_42914 <= lhs_57_fu_35642_p3;
        lhs_58_reg_42920 <= lhs_58_fu_35744_p3;
        lhs_59_reg_42926 <= lhs_59_fu_35846_p3;
        lhs_60_reg_42932 <= lhs_60_fu_35948_p3;
        lhs_61_reg_42938 <= lhs_61_fu_36050_p3;
        lhs_62_reg_42944 <= lhs_62_fu_36152_p3;
        lhs_9_reg_41674 <= lhs_9_fu_23514_p3;
        or_ln346_10_reg_40609 <= or_ln346_10_fu_17363_p2;
        or_ln346_11_reg_40624 <= or_ln346_11_fu_17507_p2;
        or_ln346_14_reg_40697 <= or_ln346_14_fu_17735_p2;
        or_ln346_18_reg_41053 <= or_ln346_18_fu_20438_p2;
        or_ln346_19_reg_41068 <= or_ln346_19_fu_20567_p2;
        or_ln346_21_reg_41083 <= or_ln346_21_fu_20845_p2;
        or_ln346_22_reg_41098 <= or_ln346_22_fu_20974_p2;
        or_ln346_23_reg_41113 <= or_ln346_23_fu_21103_p2;
        or_ln346_24_reg_40975 <= or_ln346_24_fu_18373_p2;
        or_ln346_25_reg_41128 <= or_ln346_25_fu_21249_p2;
        or_ln346_26_reg_41143 <= or_ln346_26_fu_21378_p2;
        or_ln346_2_reg_40395 <= or_ln346_2_fu_16621_p2;
        or_ln346_39_reg_41524 <= or_ln346_39_fu_22322_p2;
        or_ln346_45_reg_41766 <= or_ln346_45_fu_27058_p2;
        or_ln346_51_reg_41936 <= or_ln346_51_fu_27592_p2;
        or_ln346_53_reg_41982 <= or_ln346_53_fu_27853_p2;
        or_ln346_61_reg_42200 <= or_ln346_61_fu_28375_p2;
        or_ln346_68_reg_42551 <= or_ln346_68_fu_33151_p2;
        or_ln346_6_reg_40503 <= or_ln346_6_fu_16999_p2;
        or_ln346_76_reg_42775 <= or_ln346_76_fu_33748_p2;
        overflow_10_reg_40604 <= overflow_10_fu_17333_p2;
        overflow_11_reg_40619 <= overflow_11_fu_17477_p2;
        overflow_14_reg_40692 <= overflow_14_fu_17705_p2;
        overflow_18_reg_41048 <= overflow_18_fu_20409_p2;
        overflow_19_reg_41063 <= overflow_19_fu_20538_p2;
        overflow_21_reg_41078 <= overflow_21_fu_20816_p2;
        overflow_22_reg_41093 <= overflow_22_fu_20945_p2;
        overflow_23_reg_41108 <= overflow_23_fu_21074_p2;
        overflow_24_reg_40970 <= overflow_24_fu_18343_p2;
        overflow_25_reg_41123 <= overflow_25_fu_21220_p2;
        overflow_26_reg_41138 <= overflow_26_fu_21349_p2;
        overflow_2_reg_40390 <= overflow_2_fu_16591_p2;
        overflow_39_reg_41519 <= overflow_39_fu_22292_p2;
        overflow_45_reg_41761 <= overflow_45_fu_27028_p2;
        overflow_51_reg_41931 <= overflow_51_fu_27562_p2;
        overflow_53_reg_41977 <= overflow_53_fu_27823_p2;
        overflow_61_reg_42195 <= overflow_61_fu_28345_p2;
        overflow_68_reg_42546 <= overflow_68_fu_33121_p2;
        overflow_6_reg_40498 <= overflow_6_fu_16969_p2;
        overflow_76_reg_42770 <= overflow_76_fu_33718_p2;
        p_Result_100_reg_41365 <= r_V_31_fu_496_p2[32'd45];
        p_Result_101_reg_41371 <= r_V_31_fu_496_p2[32'd45];
        p_Result_102_reg_41382 <= p_Val2_101_fu_21894_p2[32'd22];
        p_Result_103_reg_41396 <= r_V_32_fu_499_p2[32'd55];
        p_Result_104_reg_41402 <= r_V_32_fu_499_p2[32'd55];
        p_Result_105_reg_41413 <= p_Val2_104_fu_21954_p2[32'd31];
        p_Result_106_reg_41427 <= r_V_33_fu_527_p2[32'd50];
        p_Result_107_reg_41438 <= r_V_33_fu_527_p2[32'd50];
        p_Result_109_reg_41456 <= r_V_34_fu_509_p2[32'd43];
        p_Result_10_reg_40406 <= r_V_3_fu_510_p2[32'd44];
        p_Result_110_reg_41467 <= r_V_34_fu_509_p2[32'd43];
        p_Result_112_reg_41485 <= r_V_35_fu_476_p2[32'd41];
        p_Result_113_reg_41496 <= r_V_35_fu_476_p2[32'd41];
        p_Result_118_reg_41529 <= r_V_37_fu_494_p2[32'd42];
        p_Result_119_reg_41540 <= r_V_37_fu_494_p2[32'd42];
        p_Result_11_reg_40417 <= p_Val2_11_fu_16669_p2[32'd21];
        p_Result_121_reg_41558 <= r_V_38_fu_498_p2[32'd43];
        p_Result_122_reg_41569 <= r_V_38_fu_498_p2[32'd43];
        p_Result_124_reg_41587 <= r_V_39_fu_505_p2[32'd42];
        p_Result_125_reg_41598 <= r_V_39_fu_505_p2[32'd42];
        p_Result_127_reg_41616 <= r_V_40_fu_512_p2[32'd44];
        p_Result_128_reg_41627 <= r_V_40_fu_512_p2[32'd44];
        p_Result_12_reg_40431 <= r_V_4_fu_526_p2[32'd42];
        p_Result_130_reg_41645 <= r_V_41_fu_472_p2[32'd52];
        p_Result_131_reg_41656 <= r_V_41_fu_472_p2[32'd52];
        p_Result_136_reg_41771 <= r_V_43_fu_531_p2[32'd42];
        p_Result_137_reg_41777 <= r_V_43_fu_531_p2[32'd42];
        p_Result_138_reg_41788 <= p_Val2_137_fu_27106_p2[32'd19];
        p_Result_139_reg_41802 <= r_V_44_fu_520_p2[32'd41];
        p_Result_13_reg_40437 <= r_V_4_fu_526_p2[32'd42];
        p_Result_140_reg_41808 <= r_V_44_fu_520_p2[32'd41];
        p_Result_141_reg_41819 <= p_Val2_140_fu_27170_p2[32'd18];
        p_Result_142_reg_41833 <= r_V_45_fu_506_p2[32'd44];
        p_Result_143_reg_41839 <= r_V_45_fu_506_p2[32'd44];
        p_Result_144_reg_41850 <= p_Val2_143_fu_27234_p2[32'd21];
        p_Result_145_reg_41864 <= r_V_46_fu_530_p2[32'd43];
        p_Result_146_reg_41870 <= r_V_46_fu_530_p2[32'd43];
        p_Result_147_reg_41881 <= p_Val2_146_fu_27298_p2[32'd20];
        p_Result_148_reg_41895 <= r_V_47_fu_471_p2[32'd42];
        p_Result_149_reg_41901 <= r_V_47_fu_471_p2[32'd42];
        p_Result_14_reg_40448 <= p_Val2_14_fu_16733_p2[32'd19];
        p_Result_150_reg_41912 <= p_Val2_149_fu_27362_p2[32'd19];
        p_Result_154_reg_41941 <= r_V_49_fu_480_p2[32'd42];
        p_Result_155_reg_41947 <= r_V_49_fu_480_p2[32'd42];
        p_Result_156_reg_41958 <= p_Val2_155_fu_27640_p2[32'd19];
        p_Result_15_reg_40462 <= r_V_5_fu_500_p2[32'd42];
        p_Result_160_reg_41987 <= r_V_51_fu_491_p2[32'd42];
        p_Result_161_reg_41998 <= r_V_51_fu_491_p2[32'd42];
        p_Result_163_reg_42016 <= r_V_52_fu_523_p2[32'd41];
        p_Result_164_reg_42027 <= r_V_52_fu_523_p2[32'd41];
        p_Result_166_reg_42045 <= r_V_53_fu_534_p2[32'd43];
        p_Result_167_reg_42056 <= r_V_53_fu_534_p2[32'd43];
        p_Result_169_reg_42074 <= r_V_54_fu_493_p2[32'd44];
        p_Result_16_reg_40468 <= r_V_5_fu_500_p2[32'd42];
        p_Result_170_reg_42085 <= r_V_54_fu_493_p2[32'd44];
        p_Result_172_reg_42103 <= r_V_55_fu_540_p2[32'd44];
        p_Result_173_reg_42114 <= r_V_55_fu_540_p2[32'd44];
        p_Result_175_reg_42132 <= r_V_56_fu_549_p2[32'd43];
        p_Result_176_reg_42143 <= r_V_56_fu_549_p2[32'd43];
        p_Result_178_reg_42161 <= r_V_57_fu_504_p2[32'd44];
        p_Result_179_reg_42172 <= r_V_57_fu_504_p2[32'd44];
        p_Result_17_reg_40479 <= p_Val2_17_fu_16797_p2[32'd19];
        p_Result_184_reg_42205 <= r_V_59_fu_532_p2[32'd43];
        p_Result_185_reg_42216 <= r_V_59_fu_532_p2[32'd43];
        p_Result_187_reg_42386 <= r_V_60_fu_474_p2[32'd41];
        p_Result_188_reg_42392 <= r_V_60_fu_474_p2[32'd41];
        p_Result_189_reg_42403 <= p_Val2_188_fu_32682_p2[32'd18];
        p_Result_190_reg_42417 <= r_V_61_fu_543_p2[32'd42];
        p_Result_191_reg_42423 <= r_V_61_fu_543_p2[32'd42];
        p_Result_192_reg_42434 <= p_Val2_191_fu_32746_p2[32'd19];
        p_Result_193_reg_42448 <= r_V_62_fu_477_p2[32'd43];
        p_Result_194_reg_42454 <= r_V_62_fu_477_p2[32'd43];
        p_Result_195_reg_42465 <= p_Val2_194_fu_32810_p2[32'd20];
        p_Result_196_reg_42479 <= r_V_63_fu_545_p2[32'd41];
        p_Result_197_reg_42485 <= r_V_63_fu_545_p2[32'd41];
        p_Result_198_reg_42496 <= p_Val2_197_fu_32874_p2[32'd18];
        p_Result_199_reg_42510 <= r_V_64_fu_533_p2[32'd43];
        p_Result_1_reg_40329 <= r_V_fu_519_p2[32'd46];
        p_Result_200_reg_42516 <= r_V_64_fu_533_p2[32'd43];
        p_Result_201_reg_42527 <= p_Val2_200_fu_32938_p2[32'd20];
        p_Result_205_reg_42556 <= r_V_66_fu_511_p2[32'd42];
        p_Result_206_reg_42562 <= r_V_66_fu_511_p2[32'd42];
        p_Result_207_reg_42573 <= p_Val2_206_fu_33199_p2[32'd19];
        p_Result_208_reg_42587 <= r_V_67_fu_522_p2[32'd43];
        p_Result_209_reg_42593 <= r_V_67_fu_522_p2[32'd43];
        p_Result_210_reg_42604 <= p_Val2_209_fu_33263_p2[32'd20];
        p_Result_211_reg_42618 <= r_V_68_fu_544_p2[32'd41];
        p_Result_212_reg_42624 <= r_V_68_fu_544_p2[32'd41];
        p_Result_213_reg_42635 <= p_Val2_212_fu_33327_p2[32'd18];
        p_Result_214_reg_42649 <= r_V_69_fu_529_p2[32'd43];
        p_Result_215_reg_42660 <= r_V_69_fu_529_p2[32'd43];
        p_Result_217_reg_42678 <= r_V_70_fu_516_p2[32'd42];
        p_Result_218_reg_42689 <= r_V_70_fu_516_p2[32'd42];
        p_Result_21_reg_40508 <= r_V_7_fu_537_p2[32'd56];
        p_Result_220_reg_42707 <= r_V_71_fu_517_p2[32'd41];
        p_Result_221_reg_42718 <= r_V_71_fu_517_p2[32'd41];
        p_Result_223_reg_42736 <= r_V_72_fu_525_p2[32'd42];
        p_Result_224_reg_42747 <= r_V_72_fu_525_p2[32'd42];
        p_Result_229_reg_42780 <= r_V_74_fu_495_p2[32'd40];
        p_Result_22_reg_40514 <= r_V_7_fu_537_p2[32'd55];
        p_Result_230_reg_42791 <= r_V_74_fu_495_p2[32'd40];
        p_Result_232_reg_42809 <= r_V_75_fu_539_p2[32'd39];
        p_Result_233_reg_42820 <= r_V_75_fu_539_p2[32'd39];
        p_Result_235_reg_42838 <= r_V_76_fu_484_p2[32'd45];
        p_Result_236_reg_42849 <= r_V_76_fu_484_p2[32'd45];
        p_Result_238_reg_42867 <= r_V_77_fu_486_p2[32'd53];
        p_Result_239_reg_42878 <= r_V_77_fu_486_p2[32'd53];
        p_Result_23_reg_40525 <= p_Val2_23_fu_17043_p2[32'd31];
        p_Result_24_reg_40539 <= r_V_8_fu_514_p2[32'd44];
        p_Result_25_reg_40545 <= r_V_8_fu_514_p2[32'd44];
        p_Result_26_reg_40556 <= p_Val2_26_fu_17107_p2[32'd21];
        p_Result_27_reg_40570 <= r_V_9_fu_503_p2[32'd42];
        p_Result_281_reg_41716 <= ret_V_20_fu_24346_p2[32'd32];
        p_Result_282_reg_41729 <= p_Val2_281_fu_24360_p2[32'd31];
        p_Result_289_reg_41736 <= ret_V_24_fu_24382_p2[32'd32];
        p_Result_28_reg_40581 <= r_V_9_fu_503_p2[32'd42];
        p_Result_290_reg_41749 <= p_Val2_289_fu_24396_p2[32'd31];
        p_Result_2_reg_40340 <= p_Val2_2_fu_16325_p2[32'd23];
        p_Result_313_reg_42234 <= ret_V_36_fu_30165_p2[32'd32];
        p_Result_314_reg_42247 <= p_Val2_313_fu_30179_p2[32'd31];
        p_Result_315_reg_42254 <= ret_V_37_fu_30201_p2[32'd32];
        p_Result_316_reg_42267 <= p_Val2_315_fu_30215_p2[32'd31];
        p_Result_319_reg_42280 <= ret_V_39_fu_30339_p2[32'd32];
        p_Result_320_reg_42293 <= p_Val2_319_fu_30353_p2[32'd31];
        p_Result_321_reg_42300 <= ret_V_40_fu_30375_p2[32'd32];
        p_Result_322_reg_42313 <= p_Val2_321_fu_30389_p2[32'd31];
        p_Result_323_reg_42320 <= ret_V_41_fu_30411_p2[32'd32];
        p_Result_324_reg_42333 <= p_Val2_323_fu_30425_p2[32'd31];
        p_Result_327_reg_42346 <= ret_V_43_fu_30549_p2[32'd32];
        p_Result_328_reg_42359 <= p_Val2_327_fu_30563_p2[32'd31];
        p_Result_329_reg_42366 <= ret_V_44_fu_30585_p2[32'd32];
        p_Result_330_reg_42379 <= p_Val2_329_fu_30599_p2[32'd31];
        p_Result_35_reg_40629 <= r_V_10_fu_548_p2[32'd44];
        p_Result_36_reg_40640 <= r_V_10_fu_548_p2[32'd44];
        p_Result_38_reg_40658 <= r_V_11_fu_478_p2[32'd44];
        p_Result_39_reg_40669 <= r_V_11_fu_478_p2[32'd44];
        p_Result_3_reg_40354 <= r_V_1_fu_470_p2[32'd41];
        p_Result_43_reg_40702 <= r_V_12_fu_489_p2[32'd41];
        p_Result_44_reg_40708 <= r_V_12_fu_489_p2[32'd41];
        p_Result_45_reg_40719 <= p_Val2_44_fu_17783_p2[32'd18];
        p_Result_46_reg_40733 <= r_V_13_fu_501_p2[32'd42];
        p_Result_47_reg_40744 <= r_V_13_fu_501_p2[32'd42];
        p_Result_49_reg_40762 <= r_V_14_fu_546_p2[32'd44];
        p_Result_4_reg_40360 <= r_V_1_fu_470_p2[32'd41];
        p_Result_50_reg_40773 <= r_V_14_fu_546_p2[32'd44];
        p_Result_52_reg_40791 <= r_V_15_fu_482_p2[32'd42];
        p_Result_53_reg_40802 <= r_V_15_fu_482_p2[32'd42];
        p_Result_55_reg_40820 <= r_V_16_fu_492_p2[32'd43];
        p_Result_56_reg_40831 <= r_V_16_fu_492_p2[32'd43];
        p_Result_58_reg_40849 <= r_V_17_fu_485_p2[32'd41];
        p_Result_59_reg_40860 <= r_V_17_fu_485_p2[32'd41];
        p_Result_5_reg_40371 <= p_Val2_5_fu_16389_p2[32'd18];
        p_Result_61_reg_40878 <= r_V_18_fu_481_p2[32'd42];
        p_Result_62_reg_40889 <= r_V_18_fu_481_p2[32'd42];
        p_Result_64_reg_40907 <= r_V_19_fu_473_p2[32'd42];
        p_Result_65_reg_40918 <= r_V_19_fu_473_p2[32'd42];
        p_Result_67_reg_40936 <= r_V_20_fu_515_p2[32'd37];
        p_Result_68_reg_40947 <= r_V_20_fu_515_p2[32'd37];
        p_Result_73_reg_40980 <= r_V_22_fu_535_p2[32'd44];
        p_Result_74_reg_40991 <= r_V_22_fu_535_p2[32'd44];
        p_Result_76_reg_41009 <= r_V_23_fu_518_p2[32'd42];
        p_Result_77_reg_41020 <= r_V_23_fu_518_p2[32'd42];
        p_Result_79_reg_41148 <= r_V_24_fu_508_p2[32'd55];
        p_Result_80_reg_41154 <= r_V_24_fu_508_p2[32'd55];
        p_Result_81_reg_41165 <= p_Val2_80_fu_21446_p2[32'd31];
        p_Result_82_reg_41179 <= r_V_25_fu_497_p2[32'd43];
        p_Result_83_reg_41185 <= r_V_25_fu_497_p2[32'd43];
        p_Result_84_reg_41196 <= p_Val2_83_fu_21510_p2[32'd20];
        p_Result_85_reg_41210 <= r_V_26_fu_490_p2[32'd42];
        p_Result_86_reg_41216 <= r_V_26_fu_490_p2[32'd42];
        p_Result_87_reg_41227 <= p_Val2_86_fu_21574_p2[32'd19];
        p_Result_88_reg_41241 <= r_V_27_fu_541_p2[32'd43];
        p_Result_89_reg_41247 <= r_V_27_fu_541_p2[32'd43];
        p_Result_90_reg_41258 <= p_Val2_89_fu_21638_p2[32'd20];
        p_Result_91_reg_41272 <= r_V_28_fu_521_p2[32'd42];
        p_Result_92_reg_41278 <= r_V_28_fu_521_p2[32'd42];
        p_Result_93_reg_41289 <= p_Val2_92_fu_21702_p2[32'd19];
        p_Result_94_reg_41303 <= r_V_29_fu_538_p2[32'd40];
        p_Result_95_reg_41309 <= r_V_29_fu_538_p2[32'd40];
        p_Result_96_reg_41320 <= p_Val2_95_fu_21766_p2[32'd17];
        p_Result_97_reg_41334 <= r_V_30_fu_488_p2[32'd40];
        p_Result_98_reg_41340 <= r_V_30_fu_488_p2[32'd40];
        p_Result_99_reg_41351 <= p_Val2_98_fu_21830_p2[32'd17];
        p_Result_9_reg_40400 <= r_V_3_fu_510_p2[32'd44];
        p_Result_s_reg_40323 <= r_V_fu_519_p2[32'd46];
        p_Val2_101_reg_41377 <= p_Val2_101_fu_21894_p2;
        p_Val2_104_reg_41408 <= p_Val2_104_fu_21954_p2;
        p_Val2_106_reg_41433 <= {{r_V_33_fu_527_p2[50:24]}};
        p_Val2_109_reg_41462 <= {{r_V_34_fu_509_p2[43:24]}};
        p_Val2_112_reg_41491 <= {{r_V_35_fu_476_p2[41:24]}};
        p_Val2_116_reg_41514 <= p_Val2_116_fu_22190_p2;
        p_Val2_118_reg_41535 <= {{r_V_37_fu_494_p2[42:24]}};
        p_Val2_11_reg_40412 <= p_Val2_11_fu_16669_p2;
        p_Val2_121_reg_41564 <= {{r_V_38_fu_498_p2[43:24]}};
        p_Val2_124_reg_41593 <= {{r_V_39_fu_505_p2[42:24]}};
        p_Val2_127_reg_41622 <= {{r_V_40_fu_512_p2[44:24]}};
        p_Val2_130_reg_41651 <= {{r_V_41_fu_472_p2[52:24]}};
        p_Val2_134_reg_41756 <= p_Val2_134_fu_26926_p2;
        p_Val2_137_reg_41783 <= p_Val2_137_fu_27106_p2;
        p_Val2_140_reg_41814 <= p_Val2_140_fu_27170_p2;
        p_Val2_143_reg_41845 <= p_Val2_143_fu_27234_p2;
        p_Val2_146_reg_41876 <= p_Val2_146_fu_27298_p2;
        p_Val2_149_reg_41907 <= p_Val2_149_fu_27362_p2;
        p_Val2_14_reg_40443 <= p_Val2_14_fu_16733_p2;
        p_Val2_152_reg_41926 <= p_Val2_152_fu_27460_p2;
        p_Val2_155_reg_41953 <= p_Val2_155_fu_27640_p2;
        p_Val2_158_reg_41972 <= p_Val2_158_fu_27721_p2;
        p_Val2_160_reg_41993 <= {{r_V_51_fu_491_p2[42:24]}};
        p_Val2_163_reg_42022 <= {{r_V_52_fu_523_p2[41:24]}};
        p_Val2_166_reg_42051 <= {{r_V_53_fu_534_p2[43:24]}};
        p_Val2_169_reg_42080 <= {{r_V_54_fu_493_p2[44:24]}};
        p_Val2_172_reg_42109 <= {{r_V_55_fu_540_p2[44:24]}};
        p_Val2_175_reg_42138 <= {{r_V_56_fu_549_p2[43:24]}};
        p_Val2_178_reg_42167 <= {{r_V_57_fu_504_p2[44:24]}};
        p_Val2_17_reg_40474 <= p_Val2_17_fu_16797_p2;
        p_Val2_182_reg_42190 <= p_Val2_182_fu_28243_p2;
        p_Val2_184_reg_42211 <= {{r_V_59_fu_532_p2[43:24]}};
        p_Val2_188_reg_42398 <= p_Val2_188_fu_32682_p2;
        p_Val2_191_reg_42429 <= p_Val2_191_fu_32746_p2;
        p_Val2_194_reg_42460 <= p_Val2_194_fu_32810_p2;
        p_Val2_197_reg_42491 <= p_Val2_197_fu_32874_p2;
        p_Val2_200_reg_42522 <= p_Val2_200_fu_32938_p2;
        p_Val2_203_reg_42541 <= p_Val2_203_fu_33019_p2;
        p_Val2_206_reg_42568 <= p_Val2_206_fu_33199_p2;
        p_Val2_209_reg_42599 <= p_Val2_209_fu_33263_p2;
        p_Val2_20_reg_40493 <= p_Val2_20_fu_16867_p2;
        p_Val2_212_reg_42630 <= p_Val2_212_fu_33327_p2;
        p_Val2_214_reg_42655 <= {{r_V_69_fu_529_p2[43:24]}};
        p_Val2_217_reg_42684 <= {{r_V_70_fu_516_p2[42:24]}};
        p_Val2_220_reg_42713 <= {{r_V_71_fu_517_p2[41:24]}};
        p_Val2_223_reg_42742 <= {{r_V_72_fu_525_p2[42:24]}};
        p_Val2_227_reg_42765 <= p_Val2_227_fu_33616_p2;
        p_Val2_229_reg_42786 <= {{r_V_74_fu_495_p2[40:24]}};
        p_Val2_232_reg_42815 <= {{r_V_75_fu_539_p2[39:24]}};
        p_Val2_235_reg_42844 <= {{r_V_76_fu_484_p2[45:24]}};
        p_Val2_238_reg_42873 <= {{r_V_77_fu_486_p2[53:24]}};
        p_Val2_23_reg_40520 <= p_Val2_23_fu_17043_p2;
        p_Val2_26_reg_40551 <= p_Val2_26_fu_17107_p2;
        p_Val2_281_reg_41723 <= p_Val2_281_fu_24360_p2;
        p_Val2_289_reg_41743 <= p_Val2_289_fu_24396_p2;
        p_Val2_28_reg_40576 <= {{r_V_9_fu_503_p2[42:24]}};
        p_Val2_2_reg_40335 <= p_Val2_2_fu_16325_p2;
        p_Val2_313_reg_42241 <= p_Val2_313_fu_30179_p2;
        p_Val2_315_reg_42261 <= p_Val2_315_fu_30215_p2;
        p_Val2_319_reg_42287 <= p_Val2_319_fu_30353_p2;
        p_Val2_31_reg_40599 <= p_Val2_31_fu_17231_p2;
        p_Val2_321_reg_42307 <= p_Val2_321_fu_30389_p2;
        p_Val2_323_reg_42327 <= p_Val2_323_fu_30425_p2;
        p_Val2_327_reg_42353 <= p_Val2_327_fu_30563_p2;
        p_Val2_329_reg_42373 <= p_Val2_329_fu_30599_p2;
        p_Val2_33_reg_40614 <= p_Val2_33_fu_17403_p2;
        p_Val2_35_reg_40635 <= {{r_V_10_fu_548_p2[44:24]}};
        p_Val2_38_reg_40664 <= {{r_V_11_fu_478_p2[44:24]}};
        p_Val2_41_reg_40687 <= p_Val2_41_fu_17631_p2;
        p_Val2_44_reg_40714 <= p_Val2_44_fu_17783_p2;
        p_Val2_46_reg_40739 <= {{r_V_13_fu_501_p2[42:24]}};
        p_Val2_49_reg_40768 <= {{r_V_14_fu_546_p2[44:24]}};
        p_Val2_52_reg_40797 <= {{r_V_15_fu_482_p2[42:24]}};
        p_Val2_53_reg_41043 <= p_Val2_53_fu_20321_p2;
        p_Val2_55_reg_40826 <= {{r_V_16_fu_492_p2[43:24]}};
        p_Val2_56_reg_41058 <= p_Val2_56_fu_20450_p2;
        p_Val2_58_reg_40855 <= {{r_V_17_fu_485_p2[41:24]}};
        p_Val2_5_reg_40366 <= p_Val2_5_fu_16389_p2;
        p_Val2_61_reg_40884 <= {{r_V_18_fu_481_p2[42:24]}};
        p_Val2_62_reg_41073 <= p_Val2_62_fu_20728_p2;
        p_Val2_64_reg_40913 <= {{r_V_19_fu_473_p2[42:24]}};
        p_Val2_65_reg_41088 <= p_Val2_65_fu_20857_p2;
        p_Val2_67_reg_40942 <= {{r_V_20_fu_515_p2[37:24]}};
        p_Val2_68_reg_41103 <= p_Val2_68_fu_20986_p2;
        p_Val2_71_reg_40965 <= p_Val2_71_fu_18241_p2;
        p_Val2_73_reg_40986 <= {{r_V_22_fu_535_p2[44:24]}};
        p_Val2_74_reg_41118 <= p_Val2_74_fu_21132_p2;
        p_Val2_76_reg_41015 <= {{r_V_23_fu_518_p2[42:24]}};
        p_Val2_77_reg_41133 <= p_Val2_77_fu_21261_p2;
        p_Val2_80_reg_41160 <= p_Val2_80_fu_21446_p2;
        p_Val2_83_reg_41191 <= p_Val2_83_fu_21510_p2;
        p_Val2_86_reg_41222 <= p_Val2_86_fu_21574_p2;
        p_Val2_89_reg_41253 <= p_Val2_89_fu_21638_p2;
        p_Val2_8_reg_40385 <= p_Val2_8_fu_16489_p2;
        p_Val2_92_reg_41284 <= p_Val2_92_fu_21702_p2;
        p_Val2_95_reg_41315 <= p_Val2_95_fu_21766_p2;
        p_Val2_98_reg_41346 <= p_Val2_98_fu_21830_p2;
        p_read_18_reg_40258 <= p_read8_int_reg;
        p_read_18_reg_40258_pp0_iter1_reg <= p_read_18_reg_40258;
        p_read_18_reg_40258_pp0_iter2_reg <= p_read_18_reg_40258_pp0_iter1_reg;
        p_read_19_reg_40271 <= p_read7_int_reg;
        p_read_19_reg_40271_pp0_iter1_reg <= p_read_19_reg_40271;
        p_read_19_reg_40271_pp0_iter2_reg <= p_read_19_reg_40271_pp0_iter1_reg;
        p_read_20_reg_40279 <= p_read6_int_reg;
        p_read_20_reg_40279_pp0_iter1_reg <= p_read_20_reg_40279;
        p_read_21_reg_40289 <= p_read5_int_reg;
        p_read_21_reg_40289_pp0_iter1_reg <= p_read_21_reg_40289;
        p_read_22_reg_40302 <= p_read4_int_reg;
        p_read_23_reg_40314 <= p_read3_int_reg;
        r_V_10_reg_7471 <= r_V_10_fu_548_p2;
        r_V_11_reg_7475 <= r_V_11_fu_478_p2;
        r_V_12_reg_7479 <= r_V_12_fu_489_p2;
        r_V_13_reg_7483 <= r_V_13_fu_501_p2;
        r_V_14_reg_7487 <= r_V_14_fu_546_p2;
        r_V_15_reg_7491 <= r_V_15_fu_482_p2;
        r_V_16_reg_7495 <= r_V_16_fu_492_p2;
        r_V_17_reg_7499 <= r_V_17_fu_485_p2;
        r_V_18_reg_7503 <= r_V_18_fu_481_p2;
        r_V_19_reg_7507 <= r_V_19_fu_473_p2;
        r_V_1_reg_7443 <= r_V_1_fu_470_p2;
        r_V_20_reg_7511 <= r_V_20_fu_515_p2;
        r_V_22_reg_7515 <= r_V_22_fu_535_p2;
        r_V_23_reg_7519 <= r_V_23_fu_518_p2;
        r_V_24_reg_11671 <= r_V_24_fu_508_p2;
        r_V_25_reg_11675 <= r_V_25_fu_497_p2;
        r_V_26_reg_11679 <= r_V_26_fu_490_p2;
        r_V_27_reg_11683 <= r_V_27_fu_541_p2;
        r_V_28_reg_11687 <= r_V_28_fu_521_p2;
        r_V_29_reg_11691 <= r_V_29_fu_538_p2;
        r_V_30_reg_11695 <= r_V_30_fu_488_p2;
        r_V_31_reg_11699 <= r_V_31_fu_496_p2;
        r_V_32_reg_11703 <= r_V_32_fu_499_p2;
        r_V_33_reg_11707 <= r_V_33_fu_527_p2;
        r_V_34_reg_11711 <= r_V_34_fu_509_p2;
        r_V_35_reg_11715 <= r_V_35_fu_476_p2;
        r_V_37_reg_11719 <= r_V_37_fu_494_p2;
        r_V_38_reg_11723 <= r_V_38_fu_498_p2;
        r_V_39_reg_11727 <= r_V_39_fu_505_p2;
        r_V_3_reg_7447 <= r_V_3_fu_510_p2;
        r_V_40_reg_11731 <= r_V_40_fu_512_p2;
        r_V_41_reg_11735 <= r_V_41_fu_472_p2;
        r_V_43_reg_14203 <= r_V_43_fu_531_p2;
        r_V_44_reg_14207 <= r_V_44_fu_520_p2;
        r_V_45_reg_14211 <= r_V_45_fu_506_p2;
        r_V_46_reg_14215 <= r_V_46_fu_530_p2;
        r_V_47_reg_14219 <= r_V_47_fu_471_p2;
        r_V_49_reg_14223 <= r_V_49_fu_480_p2;
        r_V_4_reg_7451 <= r_V_4_fu_526_p2;
        r_V_51_reg_14227 <= r_V_51_fu_491_p2;
        r_V_52_reg_14231 <= r_V_52_fu_523_p2;
        r_V_53_reg_14235 <= r_V_53_fu_534_p2;
        r_V_54_reg_14239 <= r_V_54_fu_493_p2;
        r_V_55_reg_14243 <= r_V_55_fu_540_p2;
        r_V_56_reg_14247 <= r_V_56_fu_549_p2;
        r_V_57_reg_14251 <= r_V_57_fu_504_p2;
        r_V_59_reg_14255 <= r_V_59_fu_532_p2;
        r_V_5_reg_7455 <= r_V_5_fu_500_p2;
        r_V_60_reg_16179 <= r_V_60_fu_474_p2;
        r_V_61_reg_16183 <= r_V_61_fu_543_p2;
        r_V_62_reg_16187 <= r_V_62_fu_477_p2;
        r_V_63_reg_16191 <= r_V_63_fu_545_p2;
        r_V_64_reg_16195 <= r_V_64_fu_533_p2;
        r_V_66_reg_16199 <= r_V_66_fu_511_p2;
        r_V_67_reg_16203 <= r_V_67_fu_522_p2;
        r_V_68_reg_16207 <= r_V_68_fu_544_p2;
        r_V_69_reg_16211 <= r_V_69_fu_529_p2;
        r_V_70_reg_16215 <= r_V_70_fu_516_p2;
        r_V_71_reg_16219 <= r_V_71_fu_517_p2;
        r_V_72_reg_16223 <= r_V_72_fu_525_p2;
        r_V_74_reg_16227 <= r_V_74_fu_495_p2;
        r_V_75_reg_16231 <= r_V_75_fu_539_p2;
        r_V_76_reg_16235 <= r_V_76_fu_484_p2;
        r_V_77_reg_16239 <= r_V_77_fu_486_p2;
        r_V_7_reg_7459 <= r_V_7_fu_537_p2;
        r_V_8_reg_7463 <= r_V_8_fu_514_p2;
        r_V_9_reg_7467 <= r_V_9_fu_503_p2;
        r_V_reg_7439 <= r_V_fu_519_p2;
        tmp_102_reg_40808 <= r_V_15_fu_482_p2[32'd23];
        tmp_108_reg_40837 <= r_V_16_fu_492_p2[32'd23];
        tmp_114_reg_40866 <= r_V_17_fu_485_p2[32'd23];
        tmp_120_reg_40895 <= r_V_18_fu_481_p2[32'd23];
        tmp_126_reg_40924 <= r_V_19_fu_473_p2[32'd23];
        tmp_132_reg_40953 <= r_V_20_fu_515_p2[32'd23];
        tmp_144_reg_40997 <= r_V_22_fu_535_p2[32'd23];
        tmp_150_reg_41026 <= r_V_23_fu_518_p2[32'd23];
        tmp_210_reg_41444 <= r_V_33_fu_527_p2[32'd23];
        tmp_216_reg_41473 <= r_V_34_fu_509_p2[32'd23];
        tmp_222_reg_41502 <= r_V_35_fu_476_p2[32'd23];
        tmp_234_reg_41546 <= r_V_37_fu_494_p2[32'd23];
        tmp_240_reg_41575 <= r_V_38_fu_498_p2[32'd23];
        tmp_246_reg_41604 <= r_V_39_fu_505_p2[32'd23];
        tmp_252_reg_41633 <= r_V_40_fu_512_p2[32'd23];
        tmp_258_reg_41662 <= r_V_41_fu_472_p2[32'd23];
        tmp_264_reg_41038 <= sub_ln823_1_fu_18475_p2[32'd23];
        tmp_264_reg_41038_pp0_iter1_reg <= tmp_264_reg_41038;
        tmp_318_reg_42004 <= r_V_51_fu_491_p2[32'd23];
        tmp_324_reg_42033 <= r_V_52_fu_523_p2[32'd23];
        tmp_330_reg_42062 <= r_V_53_fu_534_p2[32'd23];
        tmp_336_reg_42091 <= r_V_54_fu_493_p2[32'd23];
        tmp_342_reg_42120 <= r_V_55_fu_540_p2[32'd23];
        tmp_348_reg_42149 <= r_V_56_fu_549_p2[32'd23];
        tmp_354_reg_42178 <= r_V_57_fu_504_p2[32'd23];
        tmp_366_reg_42222 <= r_V_59_fu_532_p2[32'd23];
        tmp_426_reg_42666 <= r_V_69_fu_529_p2[32'd23];
        tmp_432_reg_42695 <= r_V_70_fu_516_p2[32'd23];
        tmp_438_reg_42724 <= r_V_71_fu_517_p2[32'd23];
        tmp_444_reg_42753 <= r_V_72_fu_525_p2[32'd23];
        tmp_456_reg_42797 <= r_V_74_fu_495_p2[32'd23];
        tmp_462_reg_42826 <= r_V_75_fu_539_p2[32'd23];
        tmp_468_reg_42855 <= r_V_76_fu_484_p2[32'd23];
        tmp_474_reg_42884 <= r_V_77_fu_486_p2[32'd23];
        tmp_54_reg_40587 <= r_V_9_fu_503_p2[32'd23];
        tmp_69_reg_40646 <= r_V_10_fu_548_p2[32'd23];
        tmp_75_reg_40675 <= r_V_11_fu_478_p2[32'd23];
        tmp_90_reg_40750 <= r_V_13_fu_501_p2[32'd23];
        tmp_96_reg_40779 <= r_V_14_fu_546_p2[32'd23];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= select_ln302_145_fu_39380_p3;
        ap_return_1_int_reg <= select_ln302_147_fu_39482_p3;
        ap_return_2_int_reg <= select_ln302_149_fu_39584_p3;
        ap_return_3_int_reg <= select_ln302_151_fu_39686_p3;
        ap_return_4_int_reg <= select_ln302_153_fu_39788_p3;
        ap_return_5_int_reg <= select_ln302_155_fu_39890_p3;
        ap_return_6_int_reg <= select_ln302_157_fu_39992_p3;
        ap_return_7_int_reg <= select_ln302_159_fu_40094_p3;
        ap_return_8_int_reg <= select_ln302_161_fu_40196_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        p_read1_int_reg <= p_read1;
        p_read2_int_reg <= p_read2;
        p_read3_int_reg <= p_read3;
        p_read4_int_reg <= p_read4;
        p_read5_int_reg <= p_read5;
        p_read6_int_reg <= p_read6;
        p_read7_int_reg <= p_read7;
        p_read8_int_reg <= p_read8;
        p_read_int_reg <= p_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = select_ln302_145_fu_39380_p3;
    end else begin
        ap_return_0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = select_ln302_147_fu_39482_p3;
    end else begin
        ap_return_1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = select_ln302_149_fu_39584_p3;
    end else begin
        ap_return_2 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = select_ln302_151_fu_39686_p3;
    end else begin
        ap_return_3 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = select_ln302_153_fu_39788_p3;
    end else begin
        ap_return_4 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = select_ln302_155_fu_39890_p3;
    end else begin
        ap_return_5 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = select_ln302_157_fu_39992_p3;
    end else begin
        ap_return_6 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = select_ln302_159_fu_40094_p3;
    end else begin
        ap_return_7 = 'bx;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = select_ln302_161_fu_40196_p3;
    end else begin
        ap_return_8 = 'bx;
    end
end

assign Range2_all_ones_10_fu_17251_p1 = p_read1_int_reg;

assign Range2_all_ones_10_fu_17251_p3 = Range2_all_ones_10_fu_17251_p1[32'd31];

assign Range2_all_ones_22_fu_18267_p3 = r_V_21_fu_18193_p2[32'd38];

assign Range2_all_ones_2_fu_16515_p3 = r_V_2_fu_16435_p2[32'd38];

assign Range2_all_ones_37_fu_22216_p3 = r_V_36_fu_22142_p2[32'd37];

assign Range2_all_ones_43_fu_26952_p3 = r_V_42_fu_26887_p2[32'd37];

assign Range2_all_ones_49_fu_27486_p3 = r_V_48_fu_27412_p2[32'd41];

assign Range2_all_ones_51_fu_27747_p3 = r_V_50_fu_27673_p2[32'd41];

assign Range2_all_ones_59_fu_28269_p3 = r_V_58_fu_28195_p2[32'd41];

assign Range2_all_ones_66_fu_33045_p3 = r_V_65_fu_32971_p2[32'd38];

assign Range2_all_ones_6_fu_16893_p3 = r_V_6_fu_16819_p2[32'd38];

assign Range2_all_ones_74_fu_33642_p3 = r_V_73_fu_33568_p2[32'd39];

assign and_ln891_10_fu_17303_p2 = (p_Result_31_fu_17211_p3 & and_ln891_81_fu_17297_p2);

assign and_ln891_11_fu_17453_p2 = (p_Result_33_fu_17383_p3 & and_ln891_82_fu_17447_p2);

assign and_ln891_12_fu_19653_p2 = (carry_23_fu_19607_p2 & Range2_all_ones_11_reg_40651);

assign and_ln891_13_fu_19802_p2 = (carry_25_fu_19756_p2 & Range2_all_ones_12_reg_40680);

assign and_ln891_14_fu_17681_p2 = (p_Result_41_fu_17611_p3 & and_ln891_83_fu_17675_p2);

assign and_ln891_15_fu_19945_p2 = (carry_28_fu_19900_p2 & Range2_all_ones_13_reg_40726);

assign and_ln891_16_fu_20093_p2 = (carry_30_fu_20047_p2 & Range2_all_ones_14_reg_40755);

assign and_ln891_17_fu_20242_p2 = (carry_32_fu_20196_p2 & Range2_all_ones_15_reg_40784);

assign and_ln891_18_fu_20387_p2 = (carry_34_fu_20341_p2 & Range2_all_ones_16_reg_40813);

assign and_ln891_19_fu_20516_p2 = (carry_36_fu_20470_p2 & Range2_all_ones_17_reg_40842);

assign and_ln891_1_fu_18667_p2 = (carry_3_fu_18622_p2 & Range2_all_ones_1_reg_40378);

assign and_ln891_20_fu_20649_p2 = (carry_38_fu_20603_p2 & Range2_all_ones_18_reg_40871);

assign and_ln891_21_fu_20794_p2 = (carry_40_fu_20748_p2 & Range2_all_ones_19_reg_40900);

assign and_ln891_22_fu_20923_p2 = (carry_42_fu_20877_p2 & Range2_all_ones_20_reg_40929);

assign and_ln891_23_fu_21052_p2 = (carry_44_fu_21006_p2 & Range2_all_ones_21_reg_40958);

assign and_ln891_24_fu_18319_p2 = (carry_46_fu_18261_p2 & Range2_all_ones_22_fu_18267_p3);

assign and_ln891_25_fu_21198_p2 = (carry_48_fu_21152_p2 & Range2_all_ones_23_reg_41002);

assign and_ln891_26_fu_21327_p2 = (carry_50_fu_21281_p2 & Range2_all_ones_24_reg_41031);

assign and_ln891_27_fu_24579_p2 = (carry_52_fu_24534_p2 & Range2_all_ones_25_reg_41172);

assign and_ln891_28_fu_24703_p2 = (carry_54_fu_24658_p2 & Range2_all_ones_26_reg_41203);

assign and_ln891_29_fu_24828_p2 = (carry_56_fu_24783_p2 & Range2_all_ones_27_reg_41234);

assign and_ln891_2_fu_16567_p2 = (carry_5_fu_16509_p2 & Range2_all_ones_2_fu_16515_p3);

assign and_ln891_30_fu_24953_p2 = (carry_58_fu_24908_p2 & Range2_all_ones_28_reg_41265);

assign and_ln891_31_fu_25078_p2 = (carry_60_fu_25033_p2 & Range2_all_ones_29_reg_41296);

assign and_ln891_32_fu_25203_p2 = (carry_62_fu_25158_p2 & Range2_all_ones_30_reg_41327);

assign and_ln891_33_fu_25328_p2 = (carry_64_fu_25283_p2 & Range2_all_ones_31_reg_41358);

assign and_ln891_34_fu_25453_p2 = (carry_66_fu_25408_p2 & Range2_all_ones_32_reg_41389);

assign and_ln891_35_fu_25575_p2 = (carry_68_fu_25530_p2 & Range2_all_ones_33_reg_41420);

assign and_ln891_36_fu_25722_p2 = (carry_70_fu_25676_p2 & Range2_all_ones_34_reg_41449);

assign and_ln891_37_fu_25871_p2 = (carry_72_fu_25825_p2 & Range2_all_ones_35_reg_41478);

assign and_ln891_38_fu_26020_p2 = (carry_74_fu_25974_p2 & Range2_all_ones_36_reg_41507);

assign and_ln891_39_fu_22268_p2 = (carry_76_fu_22210_p2 & Range2_all_ones_37_fu_22216_p3);

assign and_ln891_3_fu_18809_p2 = (carry_7_fu_18764_p2 & Range2_all_ones_3_reg_40424);

assign and_ln891_40_fu_26186_p2 = (carry_78_fu_26140_p2 & Range2_all_ones_38_reg_41551);

assign and_ln891_41_fu_26335_p2 = (carry_80_fu_26289_p2 & Range2_all_ones_39_reg_41580);

assign and_ln891_42_fu_26484_p2 = (carry_82_fu_26438_p2 & Range2_all_ones_40_reg_41609);

assign and_ln891_43_fu_26633_p2 = (carry_84_fu_26587_p2 & Range2_all_ones_41_reg_41638);

assign and_ln891_44_fu_26782_p2 = (carry_86_fu_26736_p2 & Range2_all_ones_42_reg_41667);

assign and_ln891_45_fu_27004_p2 = (carry_88_fu_26946_p2 & Range2_all_ones_43_fu_26952_p3);

assign and_ln891_46_fu_30683_p2 = (carry_90_fu_30638_p2 & Range2_all_ones_44_reg_41795);

assign and_ln891_47_fu_30808_p2 = (carry_92_fu_30763_p2 & Range2_all_ones_45_reg_41826);

assign and_ln891_48_fu_30933_p2 = (carry_94_fu_30888_p2 & Range2_all_ones_46_reg_41857);

assign and_ln891_49_fu_31058_p2 = (carry_96_fu_31013_p2 & Range2_all_ones_47_reg_41888);

assign and_ln891_4_fu_18934_p2 = (carry_9_fu_18889_p2 & Range2_all_ones_4_reg_40455);

assign and_ln891_50_fu_31183_p2 = (carry_98_fu_31138_p2 & Range2_all_ones_48_reg_41919);

assign and_ln891_51_fu_27538_p2 = (carry_100_fu_27480_p2 & Range2_all_ones_49_fu_27486_p3);

assign and_ln891_52_fu_31325_p2 = (carry_102_fu_31280_p2 & Range2_all_ones_50_reg_41965);

assign and_ln891_53_fu_27799_p2 = (carry_104_fu_27741_p2 & Range2_all_ones_51_fu_27747_p3);

assign and_ln891_54_fu_31490_p2 = (carry_106_fu_31444_p2 & Range2_all_ones_52_reg_42009);

assign and_ln891_55_fu_31639_p2 = (carry_108_fu_31593_p2 & Range2_all_ones_53_reg_42038);

assign and_ln891_56_fu_31788_p2 = (carry_110_fu_31742_p2 & Range2_all_ones_54_reg_42067);

assign and_ln891_57_fu_31937_p2 = (carry_112_fu_31891_p2 & Range2_all_ones_55_reg_42096);

assign and_ln891_58_fu_32086_p2 = (carry_114_fu_32040_p2 & Range2_all_ones_56_reg_42125);

assign and_ln891_59_fu_32235_p2 = (carry_116_fu_32189_p2 & Range2_all_ones_57_reg_42154);

assign and_ln891_5_fu_19059_p2 = (carry_11_fu_19014_p2 & Range2_all_ones_5_reg_40486);

assign and_ln891_60_fu_32384_p2 = (carry_118_fu_32338_p2 & Range2_all_ones_58_reg_42183);

assign and_ln891_61_fu_28321_p2 = (carry_120_fu_28263_p2 & Range2_all_ones_59_fu_28269_p3);

assign and_ln891_62_fu_32550_p2 = (carry_122_fu_32504_p2 & Range2_all_ones_60_reg_42227);

assign and_ln891_63_fu_36213_p2 = (carry_124_fu_36168_p2 & Range2_all_ones_61_reg_42410);

assign and_ln891_64_fu_36338_p2 = (carry_126_fu_36293_p2 & Range2_all_ones_62_reg_42441);

assign and_ln891_65_fu_36463_p2 = (carry_128_fu_36418_p2 & Range2_all_ones_63_reg_42472);

assign and_ln891_66_fu_36588_p2 = (carry_130_fu_36543_p2 & Range2_all_ones_64_reg_42503);

assign and_ln891_67_fu_36713_p2 = (carry_132_fu_36668_p2 & Range2_all_ones_65_reg_42534);

assign and_ln891_68_fu_33097_p2 = (carry_134_fu_33039_p2 & Range2_all_ones_66_fu_33045_p3);

assign and_ln891_69_fu_36855_p2 = (carry_136_fu_36810_p2 & Range2_all_ones_67_reg_42580);

assign and_ln891_6_fu_16945_p2 = (carry_13_fu_16887_p2 & Range2_all_ones_6_fu_16893_p3);

assign and_ln891_70_fu_36980_p2 = (carry_138_fu_36935_p2 & Range2_all_ones_68_reg_42611);

assign and_ln891_71_fu_37105_p2 = (carry_140_fu_37060_p2 & Range2_all_ones_69_reg_42642);

assign and_ln891_72_fu_37253_p2 = (carry_142_fu_37207_p2 & Range2_all_ones_70_reg_42671);

assign and_ln891_73_fu_37402_p2 = (carry_144_fu_37356_p2 & Range2_all_ones_71_reg_42700);

assign and_ln891_74_fu_37551_p2 = (carry_146_fu_37505_p2 & Range2_all_ones_72_reg_42729);

assign and_ln891_75_fu_37700_p2 = (carry_148_fu_37654_p2 & Range2_all_ones_73_reg_42758);

assign and_ln891_76_fu_33694_p2 = (carry_150_fu_33636_p2 & Range2_all_ones_74_fu_33642_p3);

assign and_ln891_77_fu_37866_p2 = (carry_152_fu_37820_p2 & Range2_all_ones_75_reg_42802);

assign and_ln891_78_fu_38015_p2 = (carry_154_fu_37969_p2 & Range2_all_ones_76_reg_42831);

assign and_ln891_79_fu_38164_p2 = (carry_156_fu_38118_p2 & Range2_all_ones_77_reg_42860);

assign and_ln891_7_fu_19198_p2 = (carry_15_fu_19153_p2 & Range2_all_ones_7_reg_40532);

assign and_ln891_80_fu_38313_p2 = (carry_158_fu_38267_p2 & Range2_all_ones_78_reg_42889);

assign and_ln891_81_fu_17297_p2 = (xor_ln896_20_fu_17245_p2 & Range2_all_ones_10_fu_17251_p3);

assign and_ln891_82_fu_17447_p2 = (xor_ln896_22_fu_17417_p2 & Range2_all_ones_10_fu_17251_p3);

assign and_ln891_83_fu_17675_p2 = (xor_ln896_28_fu_17645_p2 & Range2_all_ones_10_fu_17251_p3);

assign and_ln891_8_fu_19322_p2 = (carry_17_fu_19277_p2 & Range2_all_ones_8_reg_40563);

assign and_ln891_9_fu_19470_p2 = (carry_19_fu_19424_p2 & Range2_all_ones_9_reg_40592);

assign and_ln891_fu_18542_p2 = (carry_1_fu_18497_p2 & Range2_all_ones_reg_40347);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign carry_100_fu_27480_p2 = (xor_ln896_102_fu_27474_p2 & p_Result_152_fu_27440_p3);

assign carry_102_fu_31280_p2 = (xor_ln896_104_fu_31275_p2 & p_Result_155_reg_41947);

assign carry_104_fu_27741_p2 = (xor_ln896_106_fu_27735_p2 & p_Result_158_fu_27701_p3);

assign carry_106_fu_31444_p2 = (xor_ln896_108_fu_31438_p2 & p_Result_161_reg_41998);

assign carry_108_fu_31593_p2 = (xor_ln896_110_fu_31587_p2 & p_Result_164_reg_42027);

assign carry_110_fu_31742_p2 = (xor_ln896_112_fu_31736_p2 & p_Result_167_reg_42056);

assign carry_112_fu_31891_p2 = (xor_ln896_114_fu_31885_p2 & p_Result_170_reg_42085);

assign carry_114_fu_32040_p2 = (xor_ln896_116_fu_32034_p2 & p_Result_173_reg_42114);

assign carry_116_fu_32189_p2 = (xor_ln896_118_fu_32183_p2 & p_Result_176_reg_42143);

assign carry_118_fu_32338_p2 = (xor_ln896_120_fu_32332_p2 & p_Result_179_reg_42172);

assign carry_11_fu_19014_p2 = (xor_ln896_10_fu_19009_p2 & p_Result_16_reg_40468);

assign carry_120_fu_28263_p2 = (xor_ln896_122_fu_28257_p2 & p_Result_182_fu_28223_p3);

assign carry_122_fu_32504_p2 = (xor_ln896_124_fu_32498_p2 & p_Result_185_reg_42216);

assign carry_124_fu_36168_p2 = (xor_ln896_126_fu_36163_p2 & p_Result_188_reg_42392);

assign carry_126_fu_36293_p2 = (xor_ln896_128_fu_36288_p2 & p_Result_191_reg_42423);

assign carry_128_fu_36418_p2 = (xor_ln896_130_fu_36413_p2 & p_Result_194_reg_42454);

assign carry_130_fu_36543_p2 = (xor_ln896_132_fu_36538_p2 & p_Result_197_reg_42485);

assign carry_132_fu_36668_p2 = (xor_ln896_134_fu_36663_p2 & p_Result_200_reg_42516);

assign carry_134_fu_33039_p2 = (xor_ln896_136_fu_33033_p2 & p_Result_203_fu_32999_p3);

assign carry_136_fu_36810_p2 = (xor_ln896_138_fu_36805_p2 & p_Result_206_reg_42562);

assign carry_138_fu_36935_p2 = (xor_ln896_140_fu_36930_p2 & p_Result_209_reg_42593);

assign carry_13_fu_16887_p2 = (xor_ln896_12_fu_16881_p2 & p_Result_19_fu_16847_p3);

assign carry_140_fu_37060_p2 = (xor_ln896_142_fu_37055_p2 & p_Result_212_reg_42624);

assign carry_142_fu_37207_p2 = (xor_ln896_144_fu_37201_p2 & p_Result_215_reg_42660);

assign carry_144_fu_37356_p2 = (xor_ln896_146_fu_37350_p2 & p_Result_218_reg_42689);

assign carry_146_fu_37505_p2 = (xor_ln896_148_fu_37499_p2 & p_Result_221_reg_42718);

assign carry_148_fu_37654_p2 = (xor_ln896_150_fu_37648_p2 & p_Result_224_reg_42747);

assign carry_150_fu_33636_p2 = (xor_ln896_152_fu_33630_p2 & p_Result_227_fu_33596_p3);

assign carry_152_fu_37820_p2 = (xor_ln896_154_fu_37814_p2 & p_Result_230_reg_42791);

assign carry_154_fu_37969_p2 = (xor_ln896_156_fu_37963_p2 & p_Result_233_reg_42820);

assign carry_156_fu_38118_p2 = (xor_ln896_158_fu_38112_p2 & p_Result_236_reg_42849);

assign carry_158_fu_38267_p2 = (xor_ln896_160_fu_38261_p2 & p_Result_239_reg_42878);

assign carry_15_fu_19153_p2 = (xor_ln896_14_fu_19148_p2 & p_Result_22_reg_40514);

assign carry_17_fu_19277_p2 = (xor_ln896_16_fu_19272_p2 & p_Result_25_reg_40545);

assign carry_19_fu_19424_p2 = (xor_ln896_18_fu_19418_p2 & p_Result_28_reg_40581);

assign carry_1_fu_18497_p2 = (xor_ln896_fu_18492_p2 & p_Result_1_reg_40329);

assign carry_23_fu_19607_p2 = (xor_ln896_24_fu_19601_p2 & p_Result_36_reg_40640);

assign carry_25_fu_19756_p2 = (xor_ln896_26_fu_19750_p2 & p_Result_39_reg_40669);

assign carry_28_fu_19900_p2 = (xor_ln896_30_fu_19895_p2 & p_Result_44_reg_40708);

assign carry_30_fu_20047_p2 = (xor_ln896_32_fu_20041_p2 & p_Result_47_reg_40744);

assign carry_32_fu_20196_p2 = (xor_ln896_34_fu_20190_p2 & p_Result_50_reg_40773);

assign carry_34_fu_20341_p2 = (xor_ln896_36_fu_20335_p2 & p_Result_53_reg_40802);

assign carry_36_fu_20470_p2 = (xor_ln896_38_fu_20464_p2 & p_Result_56_reg_40831);

assign carry_38_fu_20603_p2 = (xor_ln896_40_fu_20597_p2 & p_Result_59_reg_40860);

assign carry_3_fu_18622_p2 = (xor_ln896_2_fu_18617_p2 & p_Result_4_reg_40360);

assign carry_40_fu_20748_p2 = (xor_ln896_42_fu_20742_p2 & p_Result_62_reg_40889);

assign carry_42_fu_20877_p2 = (xor_ln896_44_fu_20871_p2 & p_Result_65_reg_40918);

assign carry_44_fu_21006_p2 = (xor_ln896_46_fu_21000_p2 & p_Result_68_reg_40947);

assign carry_46_fu_18261_p2 = (xor_ln896_48_fu_18255_p2 & p_Result_71_fu_18221_p3);

assign carry_48_fu_21152_p2 = (xor_ln896_50_fu_21146_p2 & p_Result_74_reg_40991);

assign carry_50_fu_21281_p2 = (xor_ln896_52_fu_21275_p2 & p_Result_77_reg_41020);

assign carry_52_fu_24534_p2 = (xor_ln896_54_fu_24529_p2 & p_Result_80_reg_41154);

assign carry_54_fu_24658_p2 = (xor_ln896_56_fu_24653_p2 & p_Result_83_reg_41185);

assign carry_56_fu_24783_p2 = (xor_ln896_58_fu_24778_p2 & p_Result_86_reg_41216);

assign carry_58_fu_24908_p2 = (xor_ln896_60_fu_24903_p2 & p_Result_89_reg_41247);

assign carry_5_fu_16509_p2 = (xor_ln896_4_fu_16503_p2 & p_Result_7_fu_16469_p3);

assign carry_60_fu_25033_p2 = (xor_ln896_62_fu_25028_p2 & p_Result_92_reg_41278);

assign carry_62_fu_25158_p2 = (xor_ln896_64_fu_25153_p2 & p_Result_95_reg_41309);

assign carry_64_fu_25283_p2 = (xor_ln896_66_fu_25278_p2 & p_Result_98_reg_41340);

assign carry_66_fu_25408_p2 = (xor_ln896_68_fu_25403_p2 & p_Result_101_reg_41371);

assign carry_68_fu_25530_p2 = (xor_ln896_70_fu_25525_p2 & p_Result_104_reg_41402);

assign carry_70_fu_25676_p2 = (xor_ln896_72_fu_25670_p2 & p_Result_107_reg_41438);

assign carry_72_fu_25825_p2 = (xor_ln896_74_fu_25819_p2 & p_Result_110_reg_41467);

assign carry_74_fu_25974_p2 = (xor_ln896_76_fu_25968_p2 & p_Result_113_reg_41496);

assign carry_76_fu_22210_p2 = (xor_ln896_78_fu_22204_p2 & p_Result_116_fu_22170_p3);

assign carry_78_fu_26140_p2 = (xor_ln896_80_fu_26134_p2 & p_Result_119_reg_41540);

assign carry_7_fu_18764_p2 = (xor_ln896_6_fu_18759_p2 & p_Result_10_reg_40406);

assign carry_80_fu_26289_p2 = (xor_ln896_82_fu_26283_p2 & p_Result_122_reg_41569);

assign carry_82_fu_26438_p2 = (xor_ln896_84_fu_26432_p2 & p_Result_125_reg_41598);

assign carry_84_fu_26587_p2 = (xor_ln896_86_fu_26581_p2 & p_Result_128_reg_41627);

assign carry_86_fu_26736_p2 = (xor_ln896_88_fu_26730_p2 & p_Result_131_reg_41656);

assign carry_88_fu_26946_p2 = (xor_ln896_90_fu_26940_p2 & p_Result_134_fu_26915_p3);

assign carry_90_fu_30638_p2 = (xor_ln896_92_fu_30633_p2 & p_Result_137_reg_41777);

assign carry_92_fu_30763_p2 = (xor_ln896_94_fu_30758_p2 & p_Result_140_reg_41808);

assign carry_94_fu_30888_p2 = (xor_ln896_96_fu_30883_p2 & p_Result_143_reg_41839);

assign carry_96_fu_31013_p2 = (xor_ln896_98_fu_31008_p2 & p_Result_146_reg_41870);

assign carry_98_fu_31138_p2 = (xor_ln896_100_fu_31133_p2 & p_Result_149_reg_41901);

assign carry_9_fu_18889_p2 = (xor_ln896_8_fu_18884_p2 & p_Result_13_reg_40437);

assign deleted_ones_10_fu_17291_p2 = (or_ln890_fu_17285_p2 & Range2_all_ones_10_fu_17251_p3);

assign deleted_ones_11_fu_17441_p2 = (or_ln890_1_fu_17435_p2 & Range2_all_ones_10_fu_17251_p3);

assign deleted_ones_12_fu_19648_p2 = (or_ln890_13_fu_19642_p2 & Range2_all_ones_11_reg_40651);

assign deleted_ones_13_fu_19797_p2 = (or_ln890_14_fu_19791_p2 & Range2_all_ones_12_reg_40680);

assign deleted_ones_14_fu_17669_p2 = (or_ln890_2_fu_17663_p2 & Range2_all_ones_10_fu_17251_p3);

assign deleted_ones_15_fu_19940_p2 = (or_ln890_15_fu_19934_p2 & Range2_all_ones_13_reg_40726);

assign deleted_ones_16_fu_20088_p2 = (or_ln890_16_fu_20082_p2 & Range2_all_ones_14_reg_40755);

assign deleted_ones_17_fu_20237_p2 = (or_ln890_17_fu_20231_p2 & Range2_all_ones_15_reg_40784);

assign deleted_ones_18_fu_20382_p2 = (or_ln890_18_fu_20376_p2 & Range2_all_ones_16_reg_40813);

assign deleted_ones_19_fu_20511_p2 = (or_ln890_19_fu_20505_p2 & Range2_all_ones_17_reg_40842);

assign deleted_ones_1_fu_18662_p2 = (or_ln890_4_fu_18656_p2 & Range2_all_ones_1_reg_40378);

assign deleted_ones_20_fu_20644_p2 = (or_ln890_20_fu_20638_p2 & Range2_all_ones_18_reg_40871);

assign deleted_ones_21_fu_20789_p2 = (or_ln890_21_fu_20783_p2 & Range2_all_ones_19_reg_40900);

assign deleted_ones_22_fu_20918_p2 = (or_ln890_22_fu_20912_p2 & Range2_all_ones_20_reg_40929);

assign deleted_ones_23_fu_21047_p2 = (or_ln890_23_fu_21041_p2 & Range2_all_ones_21_reg_40958);

assign deleted_ones_24_fu_18313_p2 = (or_ln890_24_fu_18307_p2 & Range2_all_ones_22_fu_18267_p3);

assign deleted_ones_25_fu_21193_p2 = (or_ln890_25_fu_21187_p2 & Range2_all_ones_23_reg_41002);

assign deleted_ones_26_fu_21322_p2 = (or_ln890_26_fu_21316_p2 & Range2_all_ones_24_reg_41031);

assign deleted_ones_27_fu_24574_p2 = (or_ln890_27_fu_24568_p2 & Range2_all_ones_25_reg_41172);

assign deleted_ones_28_fu_24698_p2 = (or_ln890_28_fu_24692_p2 & Range2_all_ones_26_reg_41203);

assign deleted_ones_29_fu_24823_p2 = (or_ln890_29_fu_24817_p2 & Range2_all_ones_27_reg_41234);

assign deleted_ones_2_fu_16561_p2 = (or_ln890_5_fu_16555_p2 & Range2_all_ones_2_fu_16515_p3);

assign deleted_ones_30_fu_24948_p2 = (or_ln890_30_fu_24942_p2 & Range2_all_ones_28_reg_41265);

assign deleted_ones_31_fu_25073_p2 = (or_ln890_31_fu_25067_p2 & Range2_all_ones_29_reg_41296);

assign deleted_ones_32_fu_25198_p2 = (or_ln890_32_fu_25192_p2 & Range2_all_ones_30_reg_41327);

assign deleted_ones_33_fu_25323_p2 = (or_ln890_33_fu_25317_p2 & Range2_all_ones_31_reg_41358);

assign deleted_ones_34_fu_25448_p2 = (or_ln890_34_fu_25442_p2 & Range2_all_ones_32_reg_41389);

assign deleted_ones_35_fu_25570_p2 = (or_ln890_35_fu_25564_p2 & Range2_all_ones_33_reg_41420);

assign deleted_ones_36_fu_25717_p2 = (or_ln890_36_fu_25711_p2 & Range2_all_ones_34_reg_41449);

assign deleted_ones_37_fu_25866_p2 = (or_ln890_37_fu_25860_p2 & Range2_all_ones_35_reg_41478);

assign deleted_ones_38_fu_26015_p2 = (or_ln890_38_fu_26009_p2 & Range2_all_ones_36_reg_41507);

assign deleted_ones_39_fu_22262_p2 = (or_ln890_39_fu_22256_p2 & Range2_all_ones_37_fu_22216_p3);

assign deleted_ones_3_fu_18804_p2 = (or_ln890_6_fu_18798_p2 & Range2_all_ones_3_reg_40424);

assign deleted_ones_40_fu_26181_p2 = (or_ln890_40_fu_26175_p2 & Range2_all_ones_38_reg_41551);

assign deleted_ones_41_fu_26330_p2 = (or_ln890_41_fu_26324_p2 & Range2_all_ones_39_reg_41580);

assign deleted_ones_42_fu_26479_p2 = (or_ln890_42_fu_26473_p2 & Range2_all_ones_40_reg_41609);

assign deleted_ones_43_fu_26628_p2 = (or_ln890_43_fu_26622_p2 & Range2_all_ones_41_reg_41638);

assign deleted_ones_44_fu_26777_p2 = (or_ln890_44_fu_26771_p2 & Range2_all_ones_42_reg_41667);

assign deleted_ones_45_fu_26998_p2 = (or_ln890_45_fu_26992_p2 & Range2_all_ones_43_fu_26952_p3);

assign deleted_ones_46_fu_30678_p2 = (or_ln890_46_fu_30672_p2 & Range2_all_ones_44_reg_41795);

assign deleted_ones_47_fu_30803_p2 = (or_ln890_47_fu_30797_p2 & Range2_all_ones_45_reg_41826);

assign deleted_ones_48_fu_30928_p2 = (or_ln890_48_fu_30922_p2 & Range2_all_ones_46_reg_41857);

assign deleted_ones_49_fu_31053_p2 = (or_ln890_49_fu_31047_p2 & Range2_all_ones_47_reg_41888);

assign deleted_ones_4_fu_18929_p2 = (or_ln890_7_fu_18923_p2 & Range2_all_ones_4_reg_40455);

assign deleted_ones_50_fu_31178_p2 = (or_ln890_50_fu_31172_p2 & Range2_all_ones_48_reg_41919);

assign deleted_ones_51_fu_27532_p2 = (or_ln890_51_fu_27526_p2 & Range2_all_ones_49_fu_27486_p3);

assign deleted_ones_52_fu_31320_p2 = (or_ln890_52_fu_31314_p2 & Range2_all_ones_50_reg_41965);

assign deleted_ones_53_fu_27793_p2 = (or_ln890_53_fu_27787_p2 & Range2_all_ones_51_fu_27747_p3);

assign deleted_ones_54_fu_31485_p2 = (or_ln890_54_fu_31479_p2 & Range2_all_ones_52_reg_42009);

assign deleted_ones_55_fu_31634_p2 = (or_ln890_55_fu_31628_p2 & Range2_all_ones_53_reg_42038);

assign deleted_ones_56_fu_31783_p2 = (or_ln890_56_fu_31777_p2 & Range2_all_ones_54_reg_42067);

assign deleted_ones_57_fu_31932_p2 = (or_ln890_57_fu_31926_p2 & Range2_all_ones_55_reg_42096);

assign deleted_ones_58_fu_32081_p2 = (or_ln890_58_fu_32075_p2 & Range2_all_ones_56_reg_42125);

assign deleted_ones_59_fu_32230_p2 = (or_ln890_59_fu_32224_p2 & Range2_all_ones_57_reg_42154);

assign deleted_ones_5_fu_19054_p2 = (or_ln890_8_fu_19048_p2 & Range2_all_ones_5_reg_40486);

assign deleted_ones_60_fu_32379_p2 = (or_ln890_60_fu_32373_p2 & Range2_all_ones_58_reg_42183);

assign deleted_ones_61_fu_28315_p2 = (or_ln890_61_fu_28309_p2 & Range2_all_ones_59_fu_28269_p3);

assign deleted_ones_62_fu_32545_p2 = (or_ln890_62_fu_32539_p2 & Range2_all_ones_60_reg_42227);

assign deleted_ones_63_fu_36208_p2 = (or_ln890_63_fu_36202_p2 & Range2_all_ones_61_reg_42410);

assign deleted_ones_64_fu_36333_p2 = (or_ln890_64_fu_36327_p2 & Range2_all_ones_62_reg_42441);

assign deleted_ones_65_fu_36458_p2 = (or_ln890_65_fu_36452_p2 & Range2_all_ones_63_reg_42472);

assign deleted_ones_66_fu_36583_p2 = (or_ln890_66_fu_36577_p2 & Range2_all_ones_64_reg_42503);

assign deleted_ones_67_fu_36708_p2 = (or_ln890_67_fu_36702_p2 & Range2_all_ones_65_reg_42534);

assign deleted_ones_68_fu_33091_p2 = (or_ln890_68_fu_33085_p2 & Range2_all_ones_66_fu_33045_p3);

assign deleted_ones_69_fu_36850_p2 = (or_ln890_69_fu_36844_p2 & Range2_all_ones_67_reg_42580);

assign deleted_ones_6_fu_16939_p2 = (or_ln890_9_fu_16933_p2 & Range2_all_ones_6_fu_16893_p3);

assign deleted_ones_70_fu_36975_p2 = (or_ln890_70_fu_36969_p2 & Range2_all_ones_68_reg_42611);

assign deleted_ones_71_fu_37100_p2 = (or_ln890_71_fu_37094_p2 & Range2_all_ones_69_reg_42642);

assign deleted_ones_72_fu_37248_p2 = (or_ln890_72_fu_37242_p2 & Range2_all_ones_70_reg_42671);

assign deleted_ones_73_fu_37397_p2 = (or_ln890_73_fu_37391_p2 & Range2_all_ones_71_reg_42700);

assign deleted_ones_74_fu_37546_p2 = (or_ln890_74_fu_37540_p2 & Range2_all_ones_72_reg_42729);

assign deleted_ones_75_fu_37695_p2 = (or_ln890_75_fu_37689_p2 & Range2_all_ones_73_reg_42758);

assign deleted_ones_76_fu_33688_p2 = (or_ln890_76_fu_33682_p2 & Range2_all_ones_74_fu_33642_p3);

assign deleted_ones_77_fu_37861_p2 = (or_ln890_77_fu_37855_p2 & Range2_all_ones_75_reg_42802);

assign deleted_ones_78_fu_38010_p2 = (or_ln890_78_fu_38004_p2 & Range2_all_ones_76_reg_42831);

assign deleted_ones_79_fu_38159_p2 = (or_ln890_79_fu_38153_p2 & Range2_all_ones_77_reg_42860);

assign deleted_ones_7_fu_19193_p2 = (or_ln890_10_fu_19187_p2 & Range2_all_ones_7_reg_40532);

assign deleted_ones_80_fu_38308_p2 = (or_ln890_80_fu_38302_p2 & Range2_all_ones_78_reg_42889);

assign deleted_ones_8_fu_19317_p2 = (or_ln890_11_fu_19311_p2 & Range2_all_ones_8_reg_40563);

assign deleted_ones_9_fu_19465_p2 = (or_ln890_12_fu_19459_p2 & Range2_all_ones_9_reg_40592);

assign deleted_ones_fu_18537_p2 = (or_ln890_3_fu_18531_p2 & Range2_all_ones_reg_40347);

assign deleted_zeros_10_fu_19623_p2 = (or_ln888_13_fu_19617_p2 ^ Range2_all_ones_11_reg_40651);

assign deleted_zeros_11_fu_19772_p2 = (or_ln888_14_fu_19766_p2 ^ Range2_all_ones_12_reg_40680);

assign deleted_zeros_12_fu_19915_p2 = (or_ln888_15_fu_19910_p2 ^ Range2_all_ones_13_reg_40726);

assign deleted_zeros_13_fu_20063_p2 = (or_ln888_16_fu_20057_p2 ^ Range2_all_ones_14_reg_40755);

assign deleted_zeros_14_fu_20212_p2 = (or_ln888_17_fu_20206_p2 ^ Range2_all_ones_15_reg_40784);

assign deleted_zeros_15_fu_20357_p2 = (or_ln888_18_fu_20351_p2 ^ Range2_all_ones_16_reg_40813);

assign deleted_zeros_16_fu_20486_p2 = (or_ln888_19_fu_20480_p2 ^ Range2_all_ones_17_reg_40842);

assign deleted_zeros_17_fu_20619_p2 = (or_ln888_20_fu_20613_p2 ^ Range2_all_ones_18_reg_40871);

assign deleted_zeros_18_fu_20764_p2 = (or_ln888_21_fu_20758_p2 ^ Range2_all_ones_19_reg_40900);

assign deleted_zeros_19_fu_20893_p2 = (or_ln888_22_fu_20887_p2 ^ Range2_all_ones_20_reg_40929);

assign deleted_zeros_1_fu_18637_p2 = (or_ln888_4_fu_18632_p2 ^ Range2_all_ones_1_reg_40378);

assign deleted_zeros_20_fu_21022_p2 = (or_ln888_23_fu_21016_p2 ^ Range2_all_ones_21_reg_40958);

assign deleted_zeros_21_fu_18287_p2 = (or_ln888_24_fu_18281_p2 ^ Range2_all_ones_22_fu_18267_p3);

assign deleted_zeros_22_fu_21168_p2 = (or_ln888_25_fu_21162_p2 ^ Range2_all_ones_23_reg_41002);

assign deleted_zeros_23_fu_21297_p2 = (or_ln888_26_fu_21291_p2 ^ Range2_all_ones_24_reg_41031);

assign deleted_zeros_24_fu_24549_p2 = (or_ln888_27_fu_24544_p2 ^ Range2_all_ones_25_reg_41172);

assign deleted_zeros_25_fu_24673_p2 = (or_ln888_28_fu_24668_p2 ^ Range2_all_ones_26_reg_41203);

assign deleted_zeros_26_fu_24798_p2 = (or_ln888_29_fu_24793_p2 ^ Range2_all_ones_27_reg_41234);

assign deleted_zeros_27_fu_24923_p2 = (or_ln888_30_fu_24918_p2 ^ Range2_all_ones_28_reg_41265);

assign deleted_zeros_28_fu_25048_p2 = (or_ln888_31_fu_25043_p2 ^ Range2_all_ones_29_reg_41296);

assign deleted_zeros_29_fu_25173_p2 = (or_ln888_32_fu_25168_p2 ^ Range2_all_ones_30_reg_41327);

assign deleted_zeros_2_fu_16535_p2 = (or_ln888_5_fu_16529_p2 ^ Range2_all_ones_2_fu_16515_p3);

assign deleted_zeros_30_fu_25298_p2 = (or_ln888_33_fu_25293_p2 ^ Range2_all_ones_31_reg_41358);

assign deleted_zeros_31_fu_25423_p2 = (or_ln888_34_fu_25418_p2 ^ Range2_all_ones_32_reg_41389);

assign deleted_zeros_32_fu_25545_p2 = (or_ln888_35_fu_25540_p2 ^ Range2_all_ones_33_reg_41420);

assign deleted_zeros_33_fu_25692_p2 = (or_ln888_36_fu_25686_p2 ^ Range2_all_ones_34_reg_41449);

assign deleted_zeros_34_fu_25841_p2 = (or_ln888_37_fu_25835_p2 ^ Range2_all_ones_35_reg_41478);

assign deleted_zeros_35_fu_25990_p2 = (or_ln888_38_fu_25984_p2 ^ Range2_all_ones_36_reg_41507);

assign deleted_zeros_36_fu_22236_p2 = (or_ln888_39_fu_22230_p2 ^ Range2_all_ones_37_fu_22216_p3);

assign deleted_zeros_37_fu_26156_p2 = (or_ln888_40_fu_26150_p2 ^ Range2_all_ones_38_reg_41551);

assign deleted_zeros_38_fu_26305_p2 = (or_ln888_41_fu_26299_p2 ^ Range2_all_ones_39_reg_41580);

assign deleted_zeros_39_fu_26454_p2 = (or_ln888_42_fu_26448_p2 ^ Range2_all_ones_40_reg_41609);

assign deleted_zeros_3_fu_18779_p2 = (or_ln888_6_fu_18774_p2 ^ Range2_all_ones_3_reg_40424);

assign deleted_zeros_40_fu_26603_p2 = (or_ln888_43_fu_26597_p2 ^ Range2_all_ones_41_reg_41638);

assign deleted_zeros_41_fu_26752_p2 = (or_ln888_44_fu_26746_p2 ^ Range2_all_ones_42_reg_41667);

assign deleted_zeros_42_fu_26972_p2 = (or_ln888_45_fu_26966_p2 ^ Range2_all_ones_43_fu_26952_p3);

assign deleted_zeros_43_fu_30653_p2 = (or_ln888_46_fu_30648_p2 ^ Range2_all_ones_44_reg_41795);

assign deleted_zeros_44_fu_30778_p2 = (or_ln888_47_fu_30773_p2 ^ Range2_all_ones_45_reg_41826);

assign deleted_zeros_45_fu_30903_p2 = (or_ln888_48_fu_30898_p2 ^ Range2_all_ones_46_reg_41857);

assign deleted_zeros_46_fu_31028_p2 = (or_ln888_49_fu_31023_p2 ^ Range2_all_ones_47_reg_41888);

assign deleted_zeros_47_fu_31153_p2 = (or_ln888_50_fu_31148_p2 ^ Range2_all_ones_48_reg_41919);

assign deleted_zeros_48_fu_27506_p2 = (or_ln888_51_fu_27500_p2 ^ Range2_all_ones_49_fu_27486_p3);

assign deleted_zeros_49_fu_31295_p2 = (or_ln888_52_fu_31290_p2 ^ Range2_all_ones_50_reg_41965);

assign deleted_zeros_4_fu_18904_p2 = (or_ln888_7_fu_18899_p2 ^ Range2_all_ones_4_reg_40455);

assign deleted_zeros_50_fu_27767_p2 = (or_ln888_53_fu_27761_p2 ^ Range2_all_ones_51_fu_27747_p3);

assign deleted_zeros_51_fu_31460_p2 = (or_ln888_54_fu_31454_p2 ^ Range2_all_ones_52_reg_42009);

assign deleted_zeros_52_fu_31609_p2 = (or_ln888_55_fu_31603_p2 ^ Range2_all_ones_53_reg_42038);

assign deleted_zeros_53_fu_31758_p2 = (or_ln888_56_fu_31752_p2 ^ Range2_all_ones_54_reg_42067);

assign deleted_zeros_54_fu_31907_p2 = (or_ln888_57_fu_31901_p2 ^ Range2_all_ones_55_reg_42096);

assign deleted_zeros_55_fu_32056_p2 = (or_ln888_58_fu_32050_p2 ^ Range2_all_ones_56_reg_42125);

assign deleted_zeros_56_fu_32205_p2 = (or_ln888_59_fu_32199_p2 ^ Range2_all_ones_57_reg_42154);

assign deleted_zeros_57_fu_32354_p2 = (or_ln888_60_fu_32348_p2 ^ Range2_all_ones_58_reg_42183);

assign deleted_zeros_58_fu_28289_p2 = (or_ln888_61_fu_28283_p2 ^ Range2_all_ones_59_fu_28269_p3);

assign deleted_zeros_59_fu_32520_p2 = (or_ln888_62_fu_32514_p2 ^ Range2_all_ones_60_reg_42227);

assign deleted_zeros_5_fu_19029_p2 = (or_ln888_8_fu_19024_p2 ^ Range2_all_ones_5_reg_40486);

assign deleted_zeros_60_fu_36183_p2 = (or_ln888_63_fu_36178_p2 ^ Range2_all_ones_61_reg_42410);

assign deleted_zeros_61_fu_36308_p2 = (or_ln888_64_fu_36303_p2 ^ Range2_all_ones_62_reg_42441);

assign deleted_zeros_62_fu_36433_p2 = (or_ln888_65_fu_36428_p2 ^ Range2_all_ones_63_reg_42472);

assign deleted_zeros_63_fu_36558_p2 = (or_ln888_66_fu_36553_p2 ^ Range2_all_ones_64_reg_42503);

assign deleted_zeros_64_fu_36683_p2 = (or_ln888_67_fu_36678_p2 ^ Range2_all_ones_65_reg_42534);

assign deleted_zeros_65_fu_33065_p2 = (or_ln888_68_fu_33059_p2 ^ Range2_all_ones_66_fu_33045_p3);

assign deleted_zeros_66_fu_36825_p2 = (or_ln888_69_fu_36820_p2 ^ Range2_all_ones_67_reg_42580);

assign deleted_zeros_67_fu_36950_p2 = (or_ln888_70_fu_36945_p2 ^ Range2_all_ones_68_reg_42611);

assign deleted_zeros_68_fu_37075_p2 = (or_ln888_71_fu_37070_p2 ^ Range2_all_ones_69_reg_42642);

assign deleted_zeros_69_fu_37223_p2 = (or_ln888_72_fu_37217_p2 ^ Range2_all_ones_70_reg_42671);

assign deleted_zeros_6_fu_16913_p2 = (or_ln888_9_fu_16907_p2 ^ Range2_all_ones_6_fu_16893_p3);

assign deleted_zeros_70_fu_37372_p2 = (or_ln888_73_fu_37366_p2 ^ Range2_all_ones_71_reg_42700);

assign deleted_zeros_71_fu_37521_p2 = (or_ln888_74_fu_37515_p2 ^ Range2_all_ones_72_reg_42729);

assign deleted_zeros_72_fu_37670_p2 = (or_ln888_75_fu_37664_p2 ^ Range2_all_ones_73_reg_42758);

assign deleted_zeros_73_fu_33662_p2 = (or_ln888_76_fu_33656_p2 ^ Range2_all_ones_74_fu_33642_p3);

assign deleted_zeros_74_fu_37836_p2 = (or_ln888_77_fu_37830_p2 ^ Range2_all_ones_75_reg_42802);

assign deleted_zeros_75_fu_37985_p2 = (or_ln888_78_fu_37979_p2 ^ Range2_all_ones_76_reg_42831);

assign deleted_zeros_76_fu_38134_p2 = (or_ln888_79_fu_38128_p2 ^ Range2_all_ones_77_reg_42860);

assign deleted_zeros_77_fu_38283_p2 = (or_ln888_80_fu_38277_p2 ^ Range2_all_ones_78_reg_42889);

assign deleted_zeros_7_fu_19168_p2 = (or_ln888_10_fu_19163_p2 ^ Range2_all_ones_7_reg_40532);

assign deleted_zeros_8_fu_19292_p2 = (or_ln888_11_fu_19287_p2 ^ Range2_all_ones_8_reg_40563);

assign deleted_zeros_9_fu_19440_p2 = (or_ln888_12_fu_19434_p2 ^ Range2_all_ones_9_reg_40592);

assign deleted_zeros_fu_18512_p2 = (or_ln888_3_fu_18507_p2 ^ Range2_all_ones_reg_40347);

assign lhs_10_fu_23616_p3 = ((or_ln302_10_fu_23594_p2[0:0] == 1'b1) ? select_ln302_20_fu_23600_p3 : select_ln350_10_fu_23608_p3);

assign lhs_11_fu_23718_p3 = ((or_ln302_11_fu_23696_p2[0:0] == 1'b1) ? select_ln302_22_fu_23702_p3 : select_ln350_11_fu_23710_p3);

assign lhs_12_fu_23820_p3 = ((or_ln302_12_fu_23798_p2[0:0] == 1'b1) ? select_ln302_24_fu_23804_p3 : select_ln350_12_fu_23812_p3);

assign lhs_13_fu_23922_p3 = ((or_ln302_13_fu_23900_p2[0:0] == 1'b1) ? select_ln302_26_fu_23906_p3 : select_ln350_13_fu_23914_p3);

assign lhs_14_fu_24024_p3 = ((or_ln302_14_fu_24002_p2[0:0] == 1'b1) ? select_ln302_28_fu_24008_p3 : select_ln350_14_fu_24016_p3);

assign lhs_15_fu_24126_p3 = ((or_ln302_15_fu_24104_p2[0:0] == 1'b1) ? select_ln302_30_fu_24110_p3 : select_ln350_15_fu_24118_p3);

assign lhs_16_fu_24228_p3 = ((or_ln302_16_fu_24206_p2[0:0] == 1'b1) ? select_ln302_32_fu_24212_p3 : select_ln350_16_fu_24220_p3);

assign lhs_17_fu_24330_p3 = ((or_ln302_17_fu_24308_p2[0:0] == 1'b1) ? select_ln302_34_fu_24314_p3 : select_ln350_17_fu_24322_p3);

assign lhs_18_fu_28515_p3 = ((or_ln302_18_fu_28493_p2[0:0] == 1'b1) ? select_ln302_36_fu_28499_p3 : select_ln350_18_fu_28507_p3);

assign lhs_19_fu_28615_p3 = ((or_ln302_19_fu_28593_p2[0:0] == 1'b1) ? select_ln302_38_fu_28599_p3 : select_ln350_19_fu_28607_p3);

assign lhs_1_fu_22726_p3 = ((or_ln302_1_fu_22704_p2[0:0] == 1'b1) ? select_ln302_2_fu_22710_p3 : select_ln350_1_fu_22718_p3);

assign lhs_20_fu_28673_p3 = ((or_ln302_20_fu_28653_p2[0:0] == 1'b1) ? select_ln302_40_fu_28659_p3 : select_ln350_20_fu_28666_p3);

assign lhs_21_fu_28773_p3 = ((or_ln302_21_fu_28751_p2[0:0] == 1'b1) ? select_ln302_42_fu_28757_p3 : select_ln350_21_fu_28765_p3);

assign lhs_22_fu_28873_p3 = ((or_ln302_22_fu_28851_p2[0:0] == 1'b1) ? select_ln302_44_fu_28857_p3 : select_ln350_22_fu_28865_p3);

assign lhs_23_fu_28973_p3 = ((or_ln302_23_fu_28951_p2[0:0] == 1'b1) ? select_ln302_46_fu_28957_p3 : select_ln350_23_fu_28965_p3);

assign lhs_24_fu_29031_p3 = ((or_ln302_24_fu_29011_p2[0:0] == 1'b1) ? select_ln302_48_fu_29017_p3 : select_ln350_24_fu_29024_p3);

assign lhs_25_fu_29131_p3 = ((or_ln302_25_fu_29109_p2[0:0] == 1'b1) ? select_ln302_50_fu_29115_p3 : select_ln350_25_fu_29123_p3);

assign lhs_26_fu_29231_p3 = ((or_ln302_26_fu_29209_p2[0:0] == 1'b1) ? select_ln302_52_fu_29215_p3 : select_ln350_26_fu_29223_p3);

assign lhs_27_fu_29333_p3 = ((or_ln302_27_fu_29311_p2[0:0] == 1'b1) ? select_ln302_54_fu_29317_p3 : select_ln350_27_fu_29325_p3);

assign lhs_28_fu_29435_p3 = ((or_ln302_28_fu_29413_p2[0:0] == 1'b1) ? select_ln302_56_fu_29419_p3 : select_ln350_28_fu_29427_p3);

assign lhs_29_fu_29537_p3 = ((or_ln302_29_fu_29515_p2[0:0] == 1'b1) ? select_ln302_58_fu_29521_p3 : select_ln350_29_fu_29529_p3);

assign lhs_2_fu_22824_p3 = ((or_ln302_2_fu_22802_p2[0:0] == 1'b1) ? select_ln302_4_fu_22808_p3 : select_ln350_2_fu_22816_p3);

assign lhs_30_fu_29639_p3 = ((or_ln302_30_fu_29617_p2[0:0] == 1'b1) ? select_ln302_60_fu_29623_p3 : select_ln350_30_fu_29631_p3);

assign lhs_31_fu_29741_p3 = ((or_ln302_31_fu_29719_p2[0:0] == 1'b1) ? select_ln302_62_fu_29725_p3 : select_ln350_31_fu_29733_p3);

assign lhs_32_fu_29843_p3 = ((or_ln302_32_fu_29821_p2[0:0] == 1'b1) ? select_ln302_64_fu_29827_p3 : select_ln350_32_fu_29835_p3);

assign lhs_33_fu_29945_p3 = ((or_ln302_33_fu_29923_p2[0:0] == 1'b1) ? select_ln302_66_fu_29929_p3 : select_ln350_33_fu_29937_p3);

assign lhs_34_fu_30047_p3 = ((or_ln302_34_fu_30025_p2[0:0] == 1'b1) ? select_ln302_68_fu_30031_p3 : select_ln350_34_fu_30039_p3);

assign lhs_35_fu_30149_p3 = ((or_ln302_35_fu_30127_p2[0:0] == 1'b1) ? select_ln302_70_fu_30133_p3 : select_ln350_35_fu_30141_p3);

assign lhs_36_fu_33972_p3 = ((or_ln302_36_fu_33952_p2[0:0] == 1'b1) ? select_ln302_72_fu_33958_p3 : select_ln350_36_fu_33965_p3);

assign lhs_37_fu_34030_p3 = ((or_ln302_37_fu_34010_p2[0:0] == 1'b1) ? select_ln302_74_fu_34016_p3 : select_ln350_37_fu_34023_p3);

assign lhs_38_fu_30323_p3 = ((or_ln302_38_fu_30301_p2[0:0] == 1'b1) ? select_ln302_76_fu_30307_p3 : select_ln350_38_fu_30315_p3);

assign lhs_39_fu_34088_p3 = ((or_ln302_39_fu_34068_p2[0:0] == 1'b1) ? select_ln302_78_fu_34074_p3 : select_ln350_39_fu_34081_p3);

assign lhs_3_fu_22922_p3 = ((or_ln302_3_fu_22900_p2[0:0] == 1'b1) ? select_ln302_6_fu_22906_p3 : select_ln350_3_fu_22914_p3);

assign lhs_40_fu_34146_p3 = ((or_ln302_40_fu_34126_p2[0:0] == 1'b1) ? select_ln302_80_fu_34132_p3 : select_ln350_40_fu_34139_p3);

assign lhs_41_fu_34204_p3 = ((or_ln302_41_fu_34184_p2[0:0] == 1'b1) ? select_ln302_82_fu_34190_p3 : select_ln350_41_fu_34197_p3);

assign lhs_42_fu_30533_p3 = ((or_ln302_42_fu_30511_p2[0:0] == 1'b1) ? select_ln302_84_fu_30517_p3 : select_ln350_42_fu_30525_p3);

assign lhs_43_fu_34262_p3 = ((or_ln302_43_fu_34242_p2[0:0] == 1'b1) ? select_ln302_86_fu_34248_p3 : select_ln350_43_fu_34255_p3);

assign lhs_44_fu_34320_p3 = ((or_ln302_44_fu_34300_p2[0:0] == 1'b1) ? select_ln302_88_fu_34306_p3 : select_ln350_44_fu_34313_p3);

assign lhs_45_fu_34422_p3 = ((or_ln302_45_fu_34400_p2[0:0] == 1'b1) ? select_ln302_90_fu_34406_p3 : select_ln350_45_fu_34414_p3);

assign lhs_46_fu_34524_p3 = ((or_ln302_46_fu_34502_p2[0:0] == 1'b1) ? select_ln302_92_fu_34508_p3 : select_ln350_46_fu_34516_p3);

assign lhs_47_fu_34624_p3 = ((or_ln302_47_fu_34602_p2[0:0] == 1'b1) ? select_ln302_94_fu_34608_p3 : select_ln350_47_fu_34616_p3);

assign lhs_48_fu_34726_p3 = ((or_ln302_48_fu_34704_p2[0:0] == 1'b1) ? select_ln302_96_fu_34710_p3 : select_ln350_48_fu_34718_p3);

assign lhs_49_fu_34828_p3 = ((or_ln302_49_fu_34806_p2[0:0] == 1'b1) ? select_ln302_98_fu_34812_p3 : select_ln350_49_fu_34820_p3);

assign lhs_4_fu_23020_p3 = ((or_ln302_4_fu_22998_p2[0:0] == 1'b1) ? select_ln302_8_fu_23004_p3 : select_ln350_4_fu_23012_p3);

assign lhs_50_fu_34930_p3 = ((or_ln302_50_fu_34908_p2[0:0] == 1'b1) ? select_ln302_100_fu_34914_p3 : select_ln350_50_fu_34922_p3);

assign lhs_51_fu_35030_p3 = ((or_ln302_51_fu_35008_p2[0:0] == 1'b1) ? select_ln302_102_fu_35014_p3 : select_ln350_51_fu_35022_p3);

assign lhs_52_fu_35132_p3 = ((or_ln302_52_fu_35110_p2[0:0] == 1'b1) ? select_ln302_104_fu_35116_p3 : select_ln350_52_fu_35124_p3);

assign lhs_53_fu_35234_p3 = ((or_ln302_53_fu_35212_p2[0:0] == 1'b1) ? select_ln302_106_fu_35218_p3 : select_ln350_53_fu_35226_p3);

assign lhs_54_fu_35336_p3 = ((or_ln302_54_fu_35314_p2[0:0] == 1'b1) ? select_ln302_108_fu_35320_p3 : select_ln350_54_fu_35328_p3);

assign lhs_55_fu_35438_p3 = ((or_ln302_55_fu_35416_p2[0:0] == 1'b1) ? select_ln302_110_fu_35422_p3 : select_ln350_55_fu_35430_p3);

assign lhs_56_fu_35540_p3 = ((or_ln302_56_fu_35518_p2[0:0] == 1'b1) ? select_ln302_112_fu_35524_p3 : select_ln350_56_fu_35532_p3);

assign lhs_57_fu_35642_p3 = ((or_ln302_57_fu_35620_p2[0:0] == 1'b1) ? select_ln302_114_fu_35626_p3 : select_ln350_57_fu_35634_p3);

assign lhs_58_fu_35744_p3 = ((or_ln302_58_fu_35722_p2[0:0] == 1'b1) ? select_ln302_116_fu_35728_p3 : select_ln350_58_fu_35736_p3);

assign lhs_59_fu_35846_p3 = ((or_ln302_59_fu_35824_p2[0:0] == 1'b1) ? select_ln302_118_fu_35830_p3 : select_ln350_59_fu_35838_p3);

assign lhs_5_fu_23118_p3 = ((or_ln302_5_fu_23096_p2[0:0] == 1'b1) ? select_ln302_10_fu_23102_p3 : select_ln350_5_fu_23110_p3);

assign lhs_60_fu_35948_p3 = ((or_ln302_60_fu_35926_p2[0:0] == 1'b1) ? select_ln302_120_fu_35932_p3 : select_ln350_60_fu_35940_p3);

assign lhs_61_fu_36050_p3 = ((or_ln302_61_fu_36028_p2[0:0] == 1'b1) ? select_ln302_122_fu_36034_p3 : select_ln350_61_fu_36042_p3);

assign lhs_62_fu_36152_p3 = ((or_ln302_62_fu_36130_p2[0:0] == 1'b1) ? select_ln302_124_fu_36136_p3 : select_ln350_62_fu_36144_p3);

assign lhs_63_fu_38478_p3 = ((or_ln302_63_fu_38456_p2[0:0] == 1'b1) ? select_ln302_126_fu_38462_p3 : select_ln350_63_fu_38470_p3);

assign lhs_64_fu_38578_p3 = ((or_ln302_64_fu_38556_p2[0:0] == 1'b1) ? select_ln302_128_fu_38562_p3 : select_ln350_64_fu_38570_p3);

assign lhs_65_fu_38678_p3 = ((or_ln302_65_fu_38656_p2[0:0] == 1'b1) ? select_ln302_130_fu_38662_p3 : select_ln350_65_fu_38670_p3);

assign lhs_66_fu_38778_p3 = ((or_ln302_66_fu_38756_p2[0:0] == 1'b1) ? select_ln302_132_fu_38762_p3 : select_ln350_66_fu_38770_p3);

assign lhs_67_fu_38878_p3 = ((or_ln302_67_fu_38856_p2[0:0] == 1'b1) ? select_ln302_134_fu_38862_p3 : select_ln350_67_fu_38870_p3);

assign lhs_68_fu_38978_p3 = ((or_ln302_68_fu_38956_p2[0:0] == 1'b1) ? select_ln302_136_fu_38962_p3 : select_ln350_68_fu_38970_p3);

assign lhs_69_fu_39078_p3 = ((or_ln302_69_fu_39056_p2[0:0] == 1'b1) ? select_ln302_138_fu_39062_p3 : select_ln350_69_fu_39070_p3);

assign lhs_6_fu_23216_p3 = ((or_ln302_6_fu_23194_p2[0:0] == 1'b1) ? select_ln302_12_fu_23200_p3 : select_ln350_6_fu_23208_p3);

assign lhs_70_fu_39178_p3 = ((or_ln302_70_fu_39156_p2[0:0] == 1'b1) ? select_ln302_140_fu_39162_p3 : select_ln350_70_fu_39170_p3);

assign lhs_71_fu_39278_p3 = ((or_ln302_71_fu_39256_p2[0:0] == 1'b1) ? select_ln302_142_fu_39262_p3 : select_ln350_71_fu_39270_p3);

assign lhs_7_fu_23314_p3 = ((or_ln302_7_fu_23292_p2[0:0] == 1'b1) ? select_ln302_14_fu_23298_p3 : select_ln350_7_fu_23306_p3);

assign lhs_8_fu_23412_p3 = ((or_ln302_8_fu_23390_p2[0:0] == 1'b1) ? select_ln302_16_fu_23396_p3 : select_ln350_8_fu_23404_p3);

assign lhs_9_fu_23514_p3 = ((or_ln302_9_fu_23492_p2[0:0] == 1'b1) ? select_ln302_18_fu_23498_p3 : select_ln350_9_fu_23506_p3);

assign lhs_fu_22628_p3 = ((or_ln302_fu_22606_p2[0:0] == 1'b1) ? select_ln302_fu_22612_p3 : select_ln350_fu_22620_p3);

assign or_ln302_10_fu_23594_p2 = (xor_ln302_21_fu_23588_p2 | overflow_91_fu_23564_p2);

assign or_ln302_11_fu_23696_p2 = (xor_ln302_23_fu_23690_p2 | overflow_92_fu_23666_p2);

assign or_ln302_12_fu_23798_p2 = (xor_ln302_25_fu_23792_p2 | overflow_93_fu_23768_p2);

assign or_ln302_13_fu_23900_p2 = (xor_ln302_27_fu_23894_p2 | overflow_94_fu_23870_p2);

assign or_ln302_14_fu_24002_p2 = (xor_ln302_29_fu_23996_p2 | overflow_95_fu_23972_p2);

assign or_ln302_15_fu_24104_p2 = (xor_ln302_31_fu_24098_p2 | overflow_96_fu_24074_p2);

assign or_ln302_16_fu_24206_p2 = (xor_ln302_33_fu_24200_p2 | overflow_97_fu_24176_p2);

assign or_ln302_17_fu_24308_p2 = (xor_ln302_35_fu_24302_p2 | overflow_98_fu_24278_p2);

assign or_ln302_18_fu_28493_p2 = (xor_ln302_37_fu_28487_p2 | overflow_99_fu_28463_p2);

assign or_ln302_19_fu_28593_p2 = (xor_ln302_39_fu_28587_p2 | overflow_100_fu_28563_p2);

assign or_ln302_1_fu_22704_p2 = (xor_ln302_3_fu_22698_p2 | overflow_82_fu_22674_p2);

assign or_ln302_20_fu_28653_p2 = (xor_ln302_41_fu_28647_p2 | overflow_101_fu_28628_p2);

assign or_ln302_21_fu_28751_p2 = (xor_ln302_43_fu_28745_p2 | overflow_102_fu_28721_p2);

assign or_ln302_22_fu_28851_p2 = (xor_ln302_45_fu_28845_p2 | overflow_103_fu_28821_p2);

assign or_ln302_23_fu_28951_p2 = (xor_ln302_47_fu_28945_p2 | overflow_104_fu_28921_p2);

assign or_ln302_24_fu_29011_p2 = (xor_ln302_49_fu_29005_p2 | overflow_105_fu_28986_p2);

assign or_ln302_25_fu_29109_p2 = (xor_ln302_51_fu_29103_p2 | overflow_106_fu_29079_p2);

assign or_ln302_26_fu_29209_p2 = (xor_ln302_53_fu_29203_p2 | overflow_107_fu_29179_p2);

assign or_ln302_27_fu_29311_p2 = (xor_ln302_55_fu_29305_p2 | overflow_108_fu_29281_p2);

assign or_ln302_28_fu_29413_p2 = (xor_ln302_57_fu_29407_p2 | overflow_109_fu_29383_p2);

assign or_ln302_29_fu_29515_p2 = (xor_ln302_59_fu_29509_p2 | overflow_110_fu_29485_p2);

assign or_ln302_2_fu_22802_p2 = (xor_ln302_5_fu_22796_p2 | overflow_83_fu_22772_p2);

assign or_ln302_30_fu_29617_p2 = (xor_ln302_61_fu_29611_p2 | overflow_111_fu_29587_p2);

assign or_ln302_31_fu_29719_p2 = (xor_ln302_63_fu_29713_p2 | overflow_112_fu_29689_p2);

assign or_ln302_32_fu_29821_p2 = (xor_ln302_65_fu_29815_p2 | overflow_113_fu_29791_p2);

assign or_ln302_33_fu_29923_p2 = (xor_ln302_67_fu_29917_p2 | overflow_114_fu_29893_p2);

assign or_ln302_34_fu_30025_p2 = (xor_ln302_69_fu_30019_p2 | overflow_115_fu_29995_p2);

assign or_ln302_35_fu_30127_p2 = (xor_ln302_71_fu_30121_p2 | overflow_116_fu_30097_p2);

assign or_ln302_36_fu_33952_p2 = (xor_ln302_73_fu_33946_p2 | overflow_117_fu_33927_p2);

assign or_ln302_37_fu_34010_p2 = (xor_ln302_75_fu_34004_p2 | overflow_118_fu_33985_p2);

assign or_ln302_38_fu_30301_p2 = (xor_ln302_77_fu_30295_p2 | overflow_119_fu_30271_p2);

assign or_ln302_39_fu_34068_p2 = (xor_ln302_79_fu_34062_p2 | overflow_120_fu_34043_p2);

assign or_ln302_3_fu_22900_p2 = (xor_ln302_7_fu_22894_p2 | overflow_84_fu_22870_p2);

assign or_ln302_40_fu_34126_p2 = (xor_ln302_81_fu_34120_p2 | overflow_121_fu_34101_p2);

assign or_ln302_41_fu_34184_p2 = (xor_ln302_83_fu_34178_p2 | overflow_122_fu_34159_p2);

assign or_ln302_42_fu_30511_p2 = (xor_ln302_85_fu_30505_p2 | overflow_123_fu_30481_p2);

assign or_ln302_43_fu_34242_p2 = (xor_ln302_87_fu_34236_p2 | overflow_124_fu_34217_p2);

assign or_ln302_44_fu_34300_p2 = (xor_ln302_89_fu_34294_p2 | overflow_125_fu_34275_p2);

assign or_ln302_45_fu_34400_p2 = (xor_ln302_91_fu_34394_p2 | overflow_126_fu_34370_p2);

assign or_ln302_46_fu_34502_p2 = (xor_ln302_93_fu_34496_p2 | overflow_127_fu_34472_p2);

assign or_ln302_47_fu_34602_p2 = (xor_ln302_95_fu_34596_p2 | overflow_128_fu_34572_p2);

assign or_ln302_48_fu_34704_p2 = (xor_ln302_97_fu_34698_p2 | overflow_129_fu_34674_p2);

assign or_ln302_49_fu_34806_p2 = (xor_ln302_99_fu_34800_p2 | overflow_130_fu_34776_p2);

assign or_ln302_4_fu_22998_p2 = (xor_ln302_9_fu_22992_p2 | overflow_85_fu_22968_p2);

assign or_ln302_50_fu_34908_p2 = (xor_ln302_101_fu_34902_p2 | overflow_131_fu_34878_p2);

assign or_ln302_51_fu_35008_p2 = (xor_ln302_103_fu_35002_p2 | overflow_132_fu_34978_p2);

assign or_ln302_52_fu_35110_p2 = (xor_ln302_105_fu_35104_p2 | overflow_133_fu_35080_p2);

assign or_ln302_53_fu_35212_p2 = (xor_ln302_107_fu_35206_p2 | overflow_134_fu_35182_p2);

assign or_ln302_54_fu_35314_p2 = (xor_ln302_109_fu_35308_p2 | overflow_135_fu_35284_p2);

assign or_ln302_55_fu_35416_p2 = (xor_ln302_111_fu_35410_p2 | overflow_136_fu_35386_p2);

assign or_ln302_56_fu_35518_p2 = (xor_ln302_113_fu_35512_p2 | overflow_137_fu_35488_p2);

assign or_ln302_57_fu_35620_p2 = (xor_ln302_115_fu_35614_p2 | overflow_138_fu_35590_p2);

assign or_ln302_58_fu_35722_p2 = (xor_ln302_117_fu_35716_p2 | overflow_139_fu_35692_p2);

assign or_ln302_59_fu_35824_p2 = (xor_ln302_119_fu_35818_p2 | overflow_140_fu_35794_p2);

assign or_ln302_5_fu_23096_p2 = (xor_ln302_11_fu_23090_p2 | overflow_86_fu_23066_p2);

assign or_ln302_60_fu_35926_p2 = (xor_ln302_121_fu_35920_p2 | overflow_141_fu_35896_p2);

assign or_ln302_61_fu_36028_p2 = (xor_ln302_123_fu_36022_p2 | overflow_142_fu_35998_p2);

assign or_ln302_62_fu_36130_p2 = (xor_ln302_125_fu_36124_p2 | overflow_143_fu_36100_p2);

assign or_ln302_63_fu_38456_p2 = (xor_ln302_127_fu_38450_p2 | overflow_144_fu_38426_p2);

assign or_ln302_64_fu_38556_p2 = (xor_ln302_129_fu_38550_p2 | overflow_145_fu_38526_p2);

assign or_ln302_65_fu_38656_p2 = (xor_ln302_131_fu_38650_p2 | overflow_146_fu_38626_p2);

assign or_ln302_66_fu_38756_p2 = (xor_ln302_133_fu_38750_p2 | overflow_147_fu_38726_p2);

assign or_ln302_67_fu_38856_p2 = (xor_ln302_135_fu_38850_p2 | overflow_148_fu_38826_p2);

assign or_ln302_68_fu_38956_p2 = (xor_ln302_137_fu_38950_p2 | overflow_149_fu_38926_p2);

assign or_ln302_69_fu_39056_p2 = (xor_ln302_139_fu_39050_p2 | overflow_150_fu_39026_p2);

assign or_ln302_6_fu_23194_p2 = (xor_ln302_13_fu_23188_p2 | overflow_87_fu_23164_p2);

assign or_ln302_70_fu_39156_p2 = (xor_ln302_141_fu_39150_p2 | overflow_151_fu_39126_p2);

assign or_ln302_71_fu_39256_p2 = (xor_ln302_143_fu_39250_p2 | overflow_152_fu_39226_p2);

assign or_ln302_72_fu_39358_p2 = (xor_ln302_145_fu_39352_p2 | overflow_153_fu_39328_p2);

assign or_ln302_73_fu_39460_p2 = (xor_ln302_147_fu_39454_p2 | overflow_154_fu_39430_p2);

assign or_ln302_74_fu_39562_p2 = (xor_ln302_149_fu_39556_p2 | overflow_155_fu_39532_p2);

assign or_ln302_75_fu_39664_p2 = (xor_ln302_151_fu_39658_p2 | overflow_156_fu_39634_p2);

assign or_ln302_76_fu_39766_p2 = (xor_ln302_153_fu_39760_p2 | overflow_157_fu_39736_p2);

assign or_ln302_77_fu_39868_p2 = (xor_ln302_155_fu_39862_p2 | overflow_158_fu_39838_p2);

assign or_ln302_78_fu_39970_p2 = (xor_ln302_157_fu_39964_p2 | overflow_159_fu_39940_p2);

assign or_ln302_79_fu_40072_p2 = (xor_ln302_159_fu_40066_p2 | overflow_160_fu_40042_p2);

assign or_ln302_7_fu_23292_p2 = (xor_ln302_15_fu_23286_p2 | overflow_88_fu_23262_p2);

assign or_ln302_80_fu_40174_p2 = (xor_ln302_161_fu_40168_p2 | overflow_161_fu_40144_p2);

assign or_ln302_8_fu_23390_p2 = (xor_ln302_17_fu_23384_p2 | overflow_89_fu_23360_p2);

assign or_ln302_9_fu_23492_p2 = (xor_ln302_19_fu_23486_p2 | overflow_90_fu_23462_p2);

assign or_ln302_fu_22606_p2 = (xor_ln302_1_fu_22600_p2 | overflow_81_fu_22576_p2);

assign or_ln346_10_fu_17363_p2 = (underflow_10_fu_17357_p2 | overflow_10_fu_17333_p2);

assign or_ln346_11_fu_17507_p2 = (underflow_11_fu_17501_p2 | overflow_11_fu_17477_p2);

assign or_ln346_12_fu_19712_p2 = (underflow_12_fu_19699_p2 | overflow_12_fu_19675_p2);

assign or_ln346_13_fu_19861_p2 = (underflow_13_fu_19848_p2 | overflow_13_fu_19824_p2);

assign or_ln346_14_fu_17735_p2 = (underflow_14_fu_17729_p2 | overflow_14_fu_17705_p2);

assign or_ln346_15_fu_20003_p2 = (underflow_15_fu_19990_p2 | overflow_15_fu_19966_p2);

assign or_ln346_16_fu_20152_p2 = (underflow_16_fu_20139_p2 | overflow_16_fu_20115_p2);

assign or_ln346_17_fu_20301_p2 = (underflow_17_fu_20288_p2 | overflow_17_fu_20264_p2);

assign or_ln346_18_fu_20438_p2 = (underflow_18_fu_20433_p2 | overflow_18_fu_20409_p2);

assign or_ln346_19_fu_20567_p2 = (underflow_19_fu_20562_p2 | overflow_19_fu_20538_p2);

assign or_ln346_1_fu_18725_p2 = (underflow_1_fu_18712_p2 | overflow_1_fu_18688_p2);

assign or_ln346_20_fu_20708_p2 = (underflow_20_fu_20695_p2 | overflow_20_fu_20671_p2);

assign or_ln346_21_fu_20845_p2 = (underflow_21_fu_20840_p2 | overflow_21_fu_20816_p2);

assign or_ln346_22_fu_20974_p2 = (underflow_22_fu_20969_p2 | overflow_22_fu_20945_p2);

assign or_ln346_23_fu_21103_p2 = (underflow_23_fu_21098_p2 | overflow_23_fu_21074_p2);

assign or_ln346_24_fu_18373_p2 = (underflow_24_fu_18367_p2 | overflow_24_fu_18343_p2);

assign or_ln346_25_fu_21249_p2 = (underflow_25_fu_21244_p2 | overflow_25_fu_21220_p2);

assign or_ln346_26_fu_21378_p2 = (underflow_26_fu_21373_p2 | overflow_26_fu_21349_p2);

assign or_ln346_27_fu_24637_p2 = (underflow_27_fu_24624_p2 | overflow_27_fu_24600_p2);

assign or_ln346_28_fu_24761_p2 = (underflow_28_fu_24748_p2 | overflow_28_fu_24724_p2);

assign or_ln346_29_fu_24886_p2 = (underflow_29_fu_24873_p2 | overflow_29_fu_24849_p2);

assign or_ln346_2_fu_16621_p2 = (underflow_2_fu_16615_p2 | overflow_2_fu_16591_p2);

assign or_ln346_30_fu_25011_p2 = (underflow_30_fu_24998_p2 | overflow_30_fu_24974_p2);

assign or_ln346_31_fu_25136_p2 = (underflow_31_fu_25123_p2 | overflow_31_fu_25099_p2);

assign or_ln346_32_fu_25261_p2 = (underflow_32_fu_25248_p2 | overflow_32_fu_25224_p2);

assign or_ln346_33_fu_25386_p2 = (underflow_33_fu_25373_p2 | overflow_33_fu_25349_p2);

assign or_ln346_34_fu_25511_p2 = (underflow_34_fu_25498_p2 | overflow_34_fu_25474_p2);

assign or_ln346_35_fu_25633_p2 = (underflow_35_fu_25620_p2 | overflow_35_fu_25596_p2);

assign or_ln346_36_fu_25781_p2 = (underflow_36_fu_25768_p2 | overflow_36_fu_25744_p2);

assign or_ln346_37_fu_25930_p2 = (underflow_37_fu_25917_p2 | overflow_37_fu_25893_p2);

assign or_ln346_38_fu_26079_p2 = (underflow_38_fu_26066_p2 | overflow_38_fu_26042_p2);

assign or_ln346_39_fu_22322_p2 = (underflow_39_fu_22316_p2 | overflow_39_fu_22292_p2);

assign or_ln346_3_fu_18867_p2 = (underflow_3_fu_18854_p2 | overflow_3_fu_18830_p2);

assign or_ln346_40_fu_26245_p2 = (underflow_40_fu_26232_p2 | overflow_40_fu_26208_p2);

assign or_ln346_41_fu_26394_p2 = (underflow_41_fu_26381_p2 | overflow_41_fu_26357_p2);

assign or_ln346_42_fu_26543_p2 = (underflow_42_fu_26530_p2 | overflow_42_fu_26506_p2);

assign or_ln346_43_fu_26692_p2 = (underflow_43_fu_26679_p2 | overflow_43_fu_26655_p2);

assign or_ln346_44_fu_26841_p2 = (underflow_44_fu_26828_p2 | overflow_44_fu_26804_p2);

assign or_ln346_45_fu_27058_p2 = (underflow_45_fu_27052_p2 | overflow_45_fu_27028_p2);

assign or_ln346_46_fu_30741_p2 = (underflow_46_fu_30728_p2 | overflow_46_fu_30704_p2);

assign or_ln346_47_fu_30866_p2 = (underflow_47_fu_30853_p2 | overflow_47_fu_30829_p2);

assign or_ln346_48_fu_30991_p2 = (underflow_48_fu_30978_p2 | overflow_48_fu_30954_p2);

assign or_ln346_49_fu_31116_p2 = (underflow_49_fu_31103_p2 | overflow_49_fu_31079_p2);

assign or_ln346_4_fu_18992_p2 = (underflow_4_fu_18979_p2 | overflow_4_fu_18955_p2);

assign or_ln346_50_fu_31241_p2 = (underflow_50_fu_31228_p2 | overflow_50_fu_31204_p2);

assign or_ln346_51_fu_27592_p2 = (underflow_51_fu_27586_p2 | overflow_51_fu_27562_p2);

assign or_ln346_52_fu_31383_p2 = (underflow_52_fu_31370_p2 | overflow_52_fu_31346_p2);

assign or_ln346_53_fu_27853_p2 = (underflow_53_fu_27847_p2 | overflow_53_fu_27823_p2);

assign or_ln346_54_fu_31549_p2 = (underflow_54_fu_31536_p2 | overflow_54_fu_31512_p2);

assign or_ln346_55_fu_31698_p2 = (underflow_55_fu_31685_p2 | overflow_55_fu_31661_p2);

assign or_ln346_56_fu_31847_p2 = (underflow_56_fu_31834_p2 | overflow_56_fu_31810_p2);

assign or_ln346_57_fu_31996_p2 = (underflow_57_fu_31983_p2 | overflow_57_fu_31959_p2);

assign or_ln346_58_fu_32145_p2 = (underflow_58_fu_32132_p2 | overflow_58_fu_32108_p2);

assign or_ln346_59_fu_32294_p2 = (underflow_59_fu_32281_p2 | overflow_59_fu_32257_p2);

assign or_ln346_5_fu_19117_p2 = (underflow_5_fu_19104_p2 | overflow_5_fu_19080_p2);

assign or_ln346_60_fu_32443_p2 = (underflow_60_fu_32430_p2 | overflow_60_fu_32406_p2);

assign or_ln346_61_fu_28375_p2 = (underflow_61_fu_28369_p2 | overflow_61_fu_28345_p2);

assign or_ln346_62_fu_32609_p2 = (underflow_62_fu_32596_p2 | overflow_62_fu_32572_p2);

assign or_ln346_63_fu_36271_p2 = (underflow_63_fu_36258_p2 | overflow_63_fu_36234_p2);

assign or_ln346_64_fu_36396_p2 = (underflow_64_fu_36383_p2 | overflow_64_fu_36359_p2);

assign or_ln346_65_fu_36521_p2 = (underflow_65_fu_36508_p2 | overflow_65_fu_36484_p2);

assign or_ln346_66_fu_36646_p2 = (underflow_66_fu_36633_p2 | overflow_66_fu_36609_p2);

assign or_ln346_67_fu_36771_p2 = (underflow_67_fu_36758_p2 | overflow_67_fu_36734_p2);

assign or_ln346_68_fu_33151_p2 = (underflow_68_fu_33145_p2 | overflow_68_fu_33121_p2);

assign or_ln346_69_fu_36913_p2 = (underflow_69_fu_36900_p2 | overflow_69_fu_36876_p2);

assign or_ln346_6_fu_16999_p2 = (underflow_6_fu_16993_p2 | overflow_6_fu_16969_p2);

assign or_ln346_70_fu_37038_p2 = (underflow_70_fu_37025_p2 | overflow_70_fu_37001_p2);

assign or_ln346_71_fu_37163_p2 = (underflow_71_fu_37150_p2 | overflow_71_fu_37126_p2);

assign or_ln346_72_fu_37312_p2 = (underflow_72_fu_37299_p2 | overflow_72_fu_37275_p2);

assign or_ln346_73_fu_37461_p2 = (underflow_73_fu_37448_p2 | overflow_73_fu_37424_p2);

assign or_ln346_74_fu_37610_p2 = (underflow_74_fu_37597_p2 | overflow_74_fu_37573_p2);

assign or_ln346_75_fu_37759_p2 = (underflow_75_fu_37746_p2 | overflow_75_fu_37722_p2);

assign or_ln346_76_fu_33748_p2 = (underflow_76_fu_33742_p2 | overflow_76_fu_33718_p2);

assign or_ln346_77_fu_37925_p2 = (underflow_77_fu_37912_p2 | overflow_77_fu_37888_p2);

assign or_ln346_78_fu_38074_p2 = (underflow_78_fu_38061_p2 | overflow_78_fu_38037_p2);

assign or_ln346_79_fu_38223_p2 = (underflow_79_fu_38210_p2 | overflow_79_fu_38186_p2);

assign or_ln346_7_fu_19256_p2 = (underflow_7_fu_19243_p2 | overflow_7_fu_19219_p2);

assign or_ln346_80_fu_38372_p2 = (underflow_80_fu_38359_p2 | overflow_80_fu_38335_p2);

assign or_ln346_8_fu_19380_p2 = (underflow_8_fu_19367_p2 | overflow_8_fu_19343_p2);

assign or_ln346_9_fu_19529_p2 = (underflow_9_fu_19516_p2 | overflow_9_fu_19492_p2);

assign or_ln346_fu_18600_p2 = (underflow_fu_18587_p2 | overflow_fu_18563_p2);

assign or_ln888_10_fu_19163_p2 = (xor_ln888_17_fu_19158_p2 | p_Result_23_reg_40525);

assign or_ln888_11_fu_19287_p2 = (xor_ln888_19_fu_19282_p2 | p_Result_26_reg_40556);

assign or_ln888_12_fu_19434_p2 = (xor_ln888_21_fu_19429_p2 | p_Result_29_fu_19410_p3);

assign or_ln888_13_fu_19617_p2 = (xor_ln888_23_fu_19612_p2 | p_Result_37_fu_19593_p3);

assign or_ln888_14_fu_19766_p2 = (xor_ln888_25_fu_19761_p2 | p_Result_40_fu_19742_p3);

assign or_ln888_15_fu_19910_p2 = (xor_ln888_27_fu_19905_p2 | p_Result_45_reg_40719);

assign or_ln888_16_fu_20057_p2 = (xor_ln888_29_fu_20052_p2 | p_Result_48_fu_20033_p3);

assign or_ln888_17_fu_20206_p2 = (xor_ln888_31_fu_20201_p2 | p_Result_51_fu_20182_p3);

assign or_ln888_18_fu_20351_p2 = (xor_ln888_33_fu_20346_p2 | p_Result_54_fu_20327_p3);

assign or_ln888_19_fu_20480_p2 = (xor_ln888_35_fu_20475_p2 | p_Result_57_fu_20456_p3);

assign or_ln888_1_fu_17429_p2 = (xor_ln888_2_fu_17423_p2 | p_Result_34_fu_17409_p3);

assign or_ln888_20_fu_20613_p2 = (xor_ln888_37_fu_20608_p2 | p_Result_60_fu_20589_p3);

assign or_ln888_21_fu_20758_p2 = (xor_ln888_39_fu_20753_p2 | p_Result_63_fu_20734_p3);

assign or_ln888_22_fu_20887_p2 = (xor_ln888_41_fu_20882_p2 | p_Result_66_fu_20863_p3);

assign or_ln888_23_fu_21016_p2 = (xor_ln888_43_fu_21011_p2 | p_Result_69_fu_20992_p3);

assign or_ln888_24_fu_18281_p2 = (xor_ln888_45_fu_18275_p2 | p_Result_72_fu_18247_p3);

assign or_ln888_25_fu_21162_p2 = (xor_ln888_47_fu_21157_p2 | p_Result_75_fu_21138_p3);

assign or_ln888_26_fu_21291_p2 = (xor_ln888_49_fu_21286_p2 | p_Result_78_fu_21267_p3);

assign or_ln888_27_fu_24544_p2 = (xor_ln888_51_fu_24539_p2 | p_Result_81_reg_41165);

assign or_ln888_28_fu_24668_p2 = (xor_ln888_53_fu_24663_p2 | p_Result_84_reg_41196);

assign or_ln888_29_fu_24793_p2 = (xor_ln888_55_fu_24788_p2 | p_Result_87_reg_41227);

assign or_ln888_2_fu_17657_p2 = (xor_ln888_4_fu_17651_p2 | p_Result_42_fu_17637_p3);

assign or_ln888_30_fu_24918_p2 = (xor_ln888_57_fu_24913_p2 | p_Result_90_reg_41258);

assign or_ln888_31_fu_25043_p2 = (xor_ln888_59_fu_25038_p2 | p_Result_93_reg_41289);

assign or_ln888_32_fu_25168_p2 = (xor_ln888_61_fu_25163_p2 | p_Result_96_reg_41320);

assign or_ln888_33_fu_25293_p2 = (xor_ln888_63_fu_25288_p2 | p_Result_99_reg_41351);

assign or_ln888_34_fu_25418_p2 = (xor_ln888_65_fu_25413_p2 | p_Result_102_reg_41382);

assign or_ln888_35_fu_25540_p2 = (xor_ln888_67_fu_25535_p2 | p_Result_105_reg_41413);

assign or_ln888_36_fu_25686_p2 = (xor_ln888_69_fu_25681_p2 | p_Result_108_fu_25662_p3);

assign or_ln888_37_fu_25835_p2 = (xor_ln888_71_fu_25830_p2 | p_Result_111_fu_25811_p3);

assign or_ln888_38_fu_25984_p2 = (xor_ln888_73_fu_25979_p2 | p_Result_114_fu_25960_p3);

assign or_ln888_39_fu_22230_p2 = (xor_ln888_75_fu_22224_p2 | p_Result_117_fu_22196_p3);

assign or_ln888_3_fu_18507_p2 = (xor_ln888_1_fu_18502_p2 | p_Result_2_reg_40340);

assign or_ln888_40_fu_26150_p2 = (xor_ln888_77_fu_26145_p2 | p_Result_120_fu_26126_p3);

assign or_ln888_41_fu_26299_p2 = (xor_ln888_79_fu_26294_p2 | p_Result_123_fu_26275_p3);

assign or_ln888_42_fu_26448_p2 = (xor_ln888_81_fu_26443_p2 | p_Result_126_fu_26424_p3);

assign or_ln888_43_fu_26597_p2 = (xor_ln888_83_fu_26592_p2 | p_Result_129_fu_26573_p3);

assign or_ln888_44_fu_26746_p2 = (xor_ln888_85_fu_26741_p2 | p_Result_132_fu_26722_p3);

assign or_ln888_45_fu_26966_p2 = (xor_ln888_87_fu_26960_p2 | p_Result_135_fu_26932_p3);

assign or_ln888_46_fu_30648_p2 = (xor_ln888_89_fu_30643_p2 | p_Result_138_reg_41788);

assign or_ln888_47_fu_30773_p2 = (xor_ln888_91_fu_30768_p2 | p_Result_141_reg_41819);

assign or_ln888_48_fu_30898_p2 = (xor_ln888_93_fu_30893_p2 | p_Result_144_reg_41850);

assign or_ln888_49_fu_31023_p2 = (xor_ln888_95_fu_31018_p2 | p_Result_147_reg_41881);

assign or_ln888_4_fu_18632_p2 = (xor_ln888_5_fu_18627_p2 | p_Result_5_reg_40371);

assign or_ln888_50_fu_31148_p2 = (xor_ln888_97_fu_31143_p2 | p_Result_150_reg_41912);

assign or_ln888_51_fu_27500_p2 = (xor_ln888_99_fu_27494_p2 | p_Result_153_fu_27466_p3);

assign or_ln888_52_fu_31290_p2 = (xor_ln888_101_fu_31285_p2 | p_Result_156_reg_41958);

assign or_ln888_53_fu_27761_p2 = (xor_ln888_103_fu_27755_p2 | p_Result_159_fu_27727_p3);

assign or_ln888_54_fu_31454_p2 = (xor_ln888_105_fu_31449_p2 | p_Result_162_fu_31430_p3);

assign or_ln888_55_fu_31603_p2 = (xor_ln888_107_fu_31598_p2 | p_Result_165_fu_31579_p3);

assign or_ln888_56_fu_31752_p2 = (xor_ln888_109_fu_31747_p2 | p_Result_168_fu_31728_p3);

assign or_ln888_57_fu_31901_p2 = (xor_ln888_111_fu_31896_p2 | p_Result_171_fu_31877_p3);

assign or_ln888_58_fu_32050_p2 = (xor_ln888_113_fu_32045_p2 | p_Result_174_fu_32026_p3);

assign or_ln888_59_fu_32199_p2 = (xor_ln888_115_fu_32194_p2 | p_Result_177_fu_32175_p3);

assign or_ln888_5_fu_16529_p2 = (xor_ln888_7_fu_16523_p2 | p_Result_8_fu_16495_p3);

assign or_ln888_60_fu_32348_p2 = (xor_ln888_117_fu_32343_p2 | p_Result_180_fu_32324_p3);

assign or_ln888_61_fu_28283_p2 = (xor_ln888_119_fu_28277_p2 | p_Result_183_fu_28249_p3);

assign or_ln888_62_fu_32514_p2 = (xor_ln888_121_fu_32509_p2 | p_Result_186_fu_32490_p3);

assign or_ln888_63_fu_36178_p2 = (xor_ln888_123_fu_36173_p2 | p_Result_189_reg_42403);

assign or_ln888_64_fu_36303_p2 = (xor_ln888_125_fu_36298_p2 | p_Result_192_reg_42434);

assign or_ln888_65_fu_36428_p2 = (xor_ln888_127_fu_36423_p2 | p_Result_195_reg_42465);

assign or_ln888_66_fu_36553_p2 = (xor_ln888_129_fu_36548_p2 | p_Result_198_reg_42496);

assign or_ln888_67_fu_36678_p2 = (xor_ln888_131_fu_36673_p2 | p_Result_201_reg_42527);

assign or_ln888_68_fu_33059_p2 = (xor_ln888_133_fu_33053_p2 | p_Result_204_fu_33025_p3);

assign or_ln888_69_fu_36820_p2 = (xor_ln888_135_fu_36815_p2 | p_Result_207_reg_42573);

assign or_ln888_6_fu_18774_p2 = (xor_ln888_9_fu_18769_p2 | p_Result_11_reg_40417);

assign or_ln888_70_fu_36945_p2 = (xor_ln888_137_fu_36940_p2 | p_Result_210_reg_42604);

assign or_ln888_71_fu_37070_p2 = (xor_ln888_139_fu_37065_p2 | p_Result_213_reg_42635);

assign or_ln888_72_fu_37217_p2 = (xor_ln888_141_fu_37212_p2 | p_Result_216_fu_37193_p3);

assign or_ln888_73_fu_37366_p2 = (xor_ln888_143_fu_37361_p2 | p_Result_219_fu_37342_p3);

assign or_ln888_74_fu_37515_p2 = (xor_ln888_145_fu_37510_p2 | p_Result_222_fu_37491_p3);

assign or_ln888_75_fu_37664_p2 = (xor_ln888_147_fu_37659_p2 | p_Result_225_fu_37640_p3);

assign or_ln888_76_fu_33656_p2 = (xor_ln888_149_fu_33650_p2 | p_Result_228_fu_33622_p3);

assign or_ln888_77_fu_37830_p2 = (xor_ln888_151_fu_37825_p2 | p_Result_231_fu_37806_p3);

assign or_ln888_78_fu_37979_p2 = (xor_ln888_153_fu_37974_p2 | p_Result_234_fu_37955_p3);

assign or_ln888_79_fu_38128_p2 = (xor_ln888_155_fu_38123_p2 | p_Result_237_fu_38104_p3);

assign or_ln888_7_fu_18899_p2 = (xor_ln888_11_fu_18894_p2 | p_Result_14_reg_40448);

assign or_ln888_80_fu_38277_p2 = (xor_ln888_157_fu_38272_p2 | p_Result_240_fu_38253_p3);

assign or_ln888_8_fu_19024_p2 = (xor_ln888_13_fu_19019_p2 | p_Result_17_reg_40479);

assign or_ln888_9_fu_16907_p2 = (xor_ln888_15_fu_16901_p2 | p_Result_20_fu_16873_p3);

assign or_ln888_fu_17265_p2 = (xor_ln888_fu_17259_p2 | p_Result_32_fu_17237_p3);

assign or_ln890_10_fu_19187_p2 = (xor_ln890_7_fu_19181_p2 | or_ln888_10_fu_19163_p2);

assign or_ln890_11_fu_19311_p2 = (xor_ln890_8_fu_19305_p2 | or_ln888_11_fu_19287_p2);

assign or_ln890_12_fu_19459_p2 = (xor_ln890_9_fu_19453_p2 | or_ln888_12_fu_19434_p2);

assign or_ln890_13_fu_19642_p2 = (xor_ln890_11_fu_19636_p2 | or_ln888_13_fu_19617_p2);

assign or_ln890_14_fu_19791_p2 = (xor_ln890_12_fu_19785_p2 | or_ln888_14_fu_19766_p2);

assign or_ln890_15_fu_19934_p2 = (xor_ln890_13_fu_19928_p2 | or_ln888_15_fu_19910_p2);

assign or_ln890_16_fu_20082_p2 = (xor_ln890_14_fu_20076_p2 | or_ln888_16_fu_20057_p2);

assign or_ln890_17_fu_20231_p2 = (xor_ln890_15_fu_20225_p2 | or_ln888_17_fu_20206_p2);

assign or_ln890_18_fu_20376_p2 = (xor_ln890_16_fu_20370_p2 | or_ln888_18_fu_20351_p2);

assign or_ln890_19_fu_20505_p2 = (xor_ln890_17_fu_20499_p2 | or_ln888_19_fu_20480_p2);

assign or_ln890_1_fu_17435_p2 = (xor_ln890_10_fu_17279_p2 | or_ln888_1_fu_17429_p2);

assign or_ln890_20_fu_20638_p2 = (xor_ln890_18_fu_20632_p2 | or_ln888_20_fu_20613_p2);

assign or_ln890_21_fu_20783_p2 = (xor_ln890_19_fu_20777_p2 | or_ln888_21_fu_20758_p2);

assign or_ln890_22_fu_20912_p2 = (xor_ln890_20_fu_20906_p2 | or_ln888_22_fu_20887_p2);

assign or_ln890_23_fu_21041_p2 = (xor_ln890_21_fu_21035_p2 | or_ln888_23_fu_21016_p2);

assign or_ln890_24_fu_18307_p2 = (xor_ln890_22_fu_18301_p2 | or_ln888_24_fu_18281_p2);

assign or_ln890_25_fu_21187_p2 = (xor_ln890_23_fu_21181_p2 | or_ln888_25_fu_21162_p2);

assign or_ln890_26_fu_21316_p2 = (xor_ln890_24_fu_21310_p2 | or_ln888_26_fu_21291_p2);

assign or_ln890_27_fu_24568_p2 = (xor_ln890_25_fu_24562_p2 | or_ln888_27_fu_24544_p2);

assign or_ln890_28_fu_24692_p2 = (xor_ln890_26_fu_24686_p2 | or_ln888_28_fu_24668_p2);

assign or_ln890_29_fu_24817_p2 = (xor_ln890_27_fu_24811_p2 | or_ln888_29_fu_24793_p2);

assign or_ln890_2_fu_17663_p2 = (xor_ln890_10_fu_17279_p2 | or_ln888_2_fu_17657_p2);

assign or_ln890_30_fu_24942_p2 = (xor_ln890_28_fu_24936_p2 | or_ln888_30_fu_24918_p2);

assign or_ln890_31_fu_25067_p2 = (xor_ln890_29_fu_25061_p2 | or_ln888_31_fu_25043_p2);

assign or_ln890_32_fu_25192_p2 = (xor_ln890_30_fu_25186_p2 | or_ln888_32_fu_25168_p2);

assign or_ln890_33_fu_25317_p2 = (xor_ln890_31_fu_25311_p2 | or_ln888_33_fu_25293_p2);

assign or_ln890_34_fu_25442_p2 = (xor_ln890_32_fu_25436_p2 | or_ln888_34_fu_25418_p2);

assign or_ln890_35_fu_25564_p2 = (xor_ln890_33_fu_25558_p2 | or_ln888_35_fu_25540_p2);

assign or_ln890_36_fu_25711_p2 = (xor_ln890_34_fu_25705_p2 | or_ln888_36_fu_25686_p2);

assign or_ln890_37_fu_25860_p2 = (xor_ln890_35_fu_25854_p2 | or_ln888_37_fu_25835_p2);

assign or_ln890_38_fu_26009_p2 = (xor_ln890_36_fu_26003_p2 | or_ln888_38_fu_25984_p2);

assign or_ln890_39_fu_22256_p2 = (xor_ln890_37_fu_22250_p2 | or_ln888_39_fu_22230_p2);

assign or_ln890_3_fu_18531_p2 = (xor_ln890_fu_18525_p2 | or_ln888_3_fu_18507_p2);

assign or_ln890_40_fu_26175_p2 = (xor_ln890_38_fu_26169_p2 | or_ln888_40_fu_26150_p2);

assign or_ln890_41_fu_26324_p2 = (xor_ln890_39_fu_26318_p2 | or_ln888_41_fu_26299_p2);

assign or_ln890_42_fu_26473_p2 = (xor_ln890_40_fu_26467_p2 | or_ln888_42_fu_26448_p2);

assign or_ln890_43_fu_26622_p2 = (xor_ln890_41_fu_26616_p2 | or_ln888_43_fu_26597_p2);

assign or_ln890_44_fu_26771_p2 = (xor_ln890_42_fu_26765_p2 | or_ln888_44_fu_26746_p2);

assign or_ln890_45_fu_26992_p2 = (xor_ln890_43_fu_26986_p2 | or_ln888_45_fu_26966_p2);

assign or_ln890_46_fu_30672_p2 = (xor_ln890_44_fu_30666_p2 | or_ln888_46_fu_30648_p2);

assign or_ln890_47_fu_30797_p2 = (xor_ln890_45_fu_30791_p2 | or_ln888_47_fu_30773_p2);

assign or_ln890_48_fu_30922_p2 = (xor_ln890_46_fu_30916_p2 | or_ln888_48_fu_30898_p2);

assign or_ln890_49_fu_31047_p2 = (xor_ln890_47_fu_31041_p2 | or_ln888_49_fu_31023_p2);

assign or_ln890_4_fu_18656_p2 = (xor_ln890_1_fu_18650_p2 | or_ln888_4_fu_18632_p2);

assign or_ln890_50_fu_31172_p2 = (xor_ln890_48_fu_31166_p2 | or_ln888_50_fu_31148_p2);

assign or_ln890_51_fu_27526_p2 = (xor_ln890_49_fu_27520_p2 | or_ln888_51_fu_27500_p2);

assign or_ln890_52_fu_31314_p2 = (xor_ln890_50_fu_31308_p2 | or_ln888_52_fu_31290_p2);

assign or_ln890_53_fu_27787_p2 = (xor_ln890_51_fu_27781_p2 | or_ln888_53_fu_27761_p2);

assign or_ln890_54_fu_31479_p2 = (xor_ln890_52_fu_31473_p2 | or_ln888_54_fu_31454_p2);

assign or_ln890_55_fu_31628_p2 = (xor_ln890_53_fu_31622_p2 | or_ln888_55_fu_31603_p2);

assign or_ln890_56_fu_31777_p2 = (xor_ln890_54_fu_31771_p2 | or_ln888_56_fu_31752_p2);

assign or_ln890_57_fu_31926_p2 = (xor_ln890_55_fu_31920_p2 | or_ln888_57_fu_31901_p2);

assign or_ln890_58_fu_32075_p2 = (xor_ln890_56_fu_32069_p2 | or_ln888_58_fu_32050_p2);

assign or_ln890_59_fu_32224_p2 = (xor_ln890_57_fu_32218_p2 | or_ln888_59_fu_32199_p2);

assign or_ln890_5_fu_16555_p2 = (xor_ln890_2_fu_16549_p2 | or_ln888_5_fu_16529_p2);

assign or_ln890_60_fu_32373_p2 = (xor_ln890_58_fu_32367_p2 | or_ln888_60_fu_32348_p2);

assign or_ln890_61_fu_28309_p2 = (xor_ln890_59_fu_28303_p2 | or_ln888_61_fu_28283_p2);

assign or_ln890_62_fu_32539_p2 = (xor_ln890_60_fu_32533_p2 | or_ln888_62_fu_32514_p2);

assign or_ln890_63_fu_36202_p2 = (xor_ln890_61_fu_36196_p2 | or_ln888_63_fu_36178_p2);

assign or_ln890_64_fu_36327_p2 = (xor_ln890_62_fu_36321_p2 | or_ln888_64_fu_36303_p2);

assign or_ln890_65_fu_36452_p2 = (xor_ln890_63_fu_36446_p2 | or_ln888_65_fu_36428_p2);

assign or_ln890_66_fu_36577_p2 = (xor_ln890_64_fu_36571_p2 | or_ln888_66_fu_36553_p2);

assign or_ln890_67_fu_36702_p2 = (xor_ln890_65_fu_36696_p2 | or_ln888_67_fu_36678_p2);

assign or_ln890_68_fu_33085_p2 = (xor_ln890_66_fu_33079_p2 | or_ln888_68_fu_33059_p2);

assign or_ln890_69_fu_36844_p2 = (xor_ln890_67_fu_36838_p2 | or_ln888_69_fu_36820_p2);

assign or_ln890_6_fu_18798_p2 = (xor_ln890_3_fu_18792_p2 | or_ln888_6_fu_18774_p2);

assign or_ln890_70_fu_36969_p2 = (xor_ln890_68_fu_36963_p2 | or_ln888_70_fu_36945_p2);

assign or_ln890_71_fu_37094_p2 = (xor_ln890_69_fu_37088_p2 | or_ln888_71_fu_37070_p2);

assign or_ln890_72_fu_37242_p2 = (xor_ln890_70_fu_37236_p2 | or_ln888_72_fu_37217_p2);

assign or_ln890_73_fu_37391_p2 = (xor_ln890_71_fu_37385_p2 | or_ln888_73_fu_37366_p2);

assign or_ln890_74_fu_37540_p2 = (xor_ln890_72_fu_37534_p2 | or_ln888_74_fu_37515_p2);

assign or_ln890_75_fu_37689_p2 = (xor_ln890_73_fu_37683_p2 | or_ln888_75_fu_37664_p2);

assign or_ln890_76_fu_33682_p2 = (xor_ln890_74_fu_33676_p2 | or_ln888_76_fu_33656_p2);

assign or_ln890_77_fu_37855_p2 = (xor_ln890_75_fu_37849_p2 | or_ln888_77_fu_37830_p2);

assign or_ln890_78_fu_38004_p2 = (xor_ln890_76_fu_37998_p2 | or_ln888_78_fu_37979_p2);

assign or_ln890_79_fu_38153_p2 = (xor_ln890_77_fu_38147_p2 | or_ln888_79_fu_38128_p2);

assign or_ln890_7_fu_18923_p2 = (xor_ln890_4_fu_18917_p2 | or_ln888_7_fu_18899_p2);

assign or_ln890_80_fu_38302_p2 = (xor_ln890_78_fu_38296_p2 | or_ln888_80_fu_38277_p2);

assign or_ln890_8_fu_19048_p2 = (xor_ln890_5_fu_19042_p2 | or_ln888_8_fu_19024_p2);

assign or_ln890_9_fu_16933_p2 = (xor_ln890_6_fu_16927_p2 | or_ln888_9_fu_16907_p2);

assign or_ln890_fu_17285_p2 = (xor_ln890_10_fu_17279_p2 | or_ln888_fu_17265_p2);

assign or_ln895_10_fu_17321_p2 = (xor_ln895_20_fu_17315_p2 | p_Result_32_fu_17237_p3);

assign or_ln895_11_fu_17471_p2 = (xor_ln895_22_fu_17465_p2 | p_Result_34_fu_17409_p3);

assign or_ln895_12_fu_19664_p2 = (xor_ln895_24_fu_19658_p2 | p_Result_37_fu_19593_p3);

assign or_ln895_13_fu_19813_p2 = (xor_ln895_26_fu_19807_p2 | p_Result_40_fu_19742_p3);

assign or_ln895_14_fu_17699_p2 = (xor_ln895_28_fu_17693_p2 | p_Result_42_fu_17637_p3);

assign or_ln895_15_fu_19956_p2 = (xor_ln895_30_fu_19950_p2 | p_Result_45_reg_40719);

assign or_ln895_16_fu_20104_p2 = (xor_ln895_32_fu_20098_p2 | p_Result_48_fu_20033_p3);

assign or_ln895_17_fu_20253_p2 = (xor_ln895_34_fu_20247_p2 | p_Result_51_fu_20182_p3);

assign or_ln895_18_fu_20398_p2 = (xor_ln895_36_fu_20392_p2 | p_Result_54_fu_20327_p3);

assign or_ln895_19_fu_20527_p2 = (xor_ln895_38_fu_20521_p2 | p_Result_57_fu_20456_p3);

assign or_ln895_1_fu_18678_p2 = (xor_ln895_2_fu_18672_p2 | p_Result_5_reg_40371);

assign or_ln895_20_fu_20660_p2 = (xor_ln895_40_fu_20654_p2 | p_Result_60_fu_20589_p3);

assign or_ln895_21_fu_20805_p2 = (xor_ln895_42_fu_20799_p2 | p_Result_63_fu_20734_p3);

assign or_ln895_22_fu_20934_p2 = (xor_ln895_44_fu_20928_p2 | p_Result_66_fu_20863_p3);

assign or_ln895_23_fu_21063_p2 = (xor_ln895_46_fu_21057_p2 | p_Result_69_fu_20992_p3);

assign or_ln895_24_fu_18331_p2 = (xor_ln895_48_fu_18325_p2 | p_Result_72_fu_18247_p3);

assign or_ln895_25_fu_21209_p2 = (xor_ln895_50_fu_21203_p2 | p_Result_75_fu_21138_p3);

assign or_ln895_26_fu_21338_p2 = (xor_ln895_52_fu_21332_p2 | p_Result_78_fu_21267_p3);

assign or_ln895_27_fu_24590_p2 = (xor_ln895_54_fu_24584_p2 | p_Result_81_reg_41165);

assign or_ln895_28_fu_24714_p2 = (xor_ln895_56_fu_24708_p2 | p_Result_84_reg_41196);

assign or_ln895_29_fu_24839_p2 = (xor_ln895_58_fu_24833_p2 | p_Result_87_reg_41227);

assign or_ln895_2_fu_16579_p2 = (xor_ln895_4_fu_16573_p2 | p_Result_8_fu_16495_p3);

assign or_ln895_30_fu_24964_p2 = (xor_ln895_60_fu_24958_p2 | p_Result_90_reg_41258);

assign or_ln895_31_fu_25089_p2 = (xor_ln895_62_fu_25083_p2 | p_Result_93_reg_41289);

assign or_ln895_32_fu_25214_p2 = (xor_ln895_64_fu_25208_p2 | p_Result_96_reg_41320);

assign or_ln895_33_fu_25339_p2 = (xor_ln895_66_fu_25333_p2 | p_Result_99_reg_41351);

assign or_ln895_34_fu_25464_p2 = (xor_ln895_68_fu_25458_p2 | p_Result_102_reg_41382);

assign or_ln895_35_fu_25586_p2 = (xor_ln895_70_fu_25580_p2 | p_Result_105_reg_41413);

assign or_ln895_36_fu_25733_p2 = (xor_ln895_72_fu_25727_p2 | p_Result_108_fu_25662_p3);

assign or_ln895_37_fu_25882_p2 = (xor_ln895_74_fu_25876_p2 | p_Result_111_fu_25811_p3);

assign or_ln895_38_fu_26031_p2 = (xor_ln895_76_fu_26025_p2 | p_Result_114_fu_25960_p3);

assign or_ln895_39_fu_22280_p2 = (xor_ln895_78_fu_22274_p2 | p_Result_117_fu_22196_p3);

assign or_ln895_3_fu_18820_p2 = (xor_ln895_6_fu_18814_p2 | p_Result_11_reg_40417);

assign or_ln895_40_fu_26197_p2 = (xor_ln895_80_fu_26191_p2 | p_Result_120_fu_26126_p3);

assign or_ln895_41_fu_26346_p2 = (xor_ln895_82_fu_26340_p2 | p_Result_123_fu_26275_p3);

assign or_ln895_42_fu_26495_p2 = (xor_ln895_84_fu_26489_p2 | p_Result_126_fu_26424_p3);

assign or_ln895_43_fu_26644_p2 = (xor_ln895_86_fu_26638_p2 | p_Result_129_fu_26573_p3);

assign or_ln895_44_fu_26793_p2 = (xor_ln895_88_fu_26787_p2 | p_Result_132_fu_26722_p3);

assign or_ln895_45_fu_27016_p2 = (xor_ln895_90_fu_27010_p2 | p_Result_135_fu_26932_p3);

assign or_ln895_46_fu_30694_p2 = (xor_ln895_92_fu_30688_p2 | p_Result_138_reg_41788);

assign or_ln895_47_fu_30819_p2 = (xor_ln895_94_fu_30813_p2 | p_Result_141_reg_41819);

assign or_ln895_48_fu_30944_p2 = (xor_ln895_96_fu_30938_p2 | p_Result_144_reg_41850);

assign or_ln895_49_fu_31069_p2 = (xor_ln895_98_fu_31063_p2 | p_Result_147_reg_41881);

assign or_ln895_4_fu_18945_p2 = (xor_ln895_8_fu_18939_p2 | p_Result_14_reg_40448);

assign or_ln895_50_fu_31194_p2 = (xor_ln895_100_fu_31188_p2 | p_Result_150_reg_41912);

assign or_ln895_51_fu_27550_p2 = (xor_ln895_102_fu_27544_p2 | p_Result_153_fu_27466_p3);

assign or_ln895_52_fu_31336_p2 = (xor_ln895_104_fu_31330_p2 | p_Result_156_reg_41958);

assign or_ln895_53_fu_27811_p2 = (xor_ln895_106_fu_27805_p2 | p_Result_159_fu_27727_p3);

assign or_ln895_54_fu_31501_p2 = (xor_ln895_108_fu_31495_p2 | p_Result_162_fu_31430_p3);

assign or_ln895_55_fu_31650_p2 = (xor_ln895_110_fu_31644_p2 | p_Result_165_fu_31579_p3);

assign or_ln895_56_fu_31799_p2 = (xor_ln895_112_fu_31793_p2 | p_Result_168_fu_31728_p3);

assign or_ln895_57_fu_31948_p2 = (xor_ln895_114_fu_31942_p2 | p_Result_171_fu_31877_p3);

assign or_ln895_58_fu_32097_p2 = (xor_ln895_116_fu_32091_p2 | p_Result_174_fu_32026_p3);

assign or_ln895_59_fu_32246_p2 = (xor_ln895_118_fu_32240_p2 | p_Result_177_fu_32175_p3);

assign or_ln895_5_fu_19070_p2 = (xor_ln895_10_fu_19064_p2 | p_Result_17_reg_40479);

assign or_ln895_60_fu_32395_p2 = (xor_ln895_120_fu_32389_p2 | p_Result_180_fu_32324_p3);

assign or_ln895_61_fu_28333_p2 = (xor_ln895_122_fu_28327_p2 | p_Result_183_fu_28249_p3);

assign or_ln895_62_fu_32561_p2 = (xor_ln895_124_fu_32555_p2 | p_Result_186_fu_32490_p3);

assign or_ln895_63_fu_36224_p2 = (xor_ln895_126_fu_36218_p2 | p_Result_189_reg_42403);

assign or_ln895_64_fu_36349_p2 = (xor_ln895_128_fu_36343_p2 | p_Result_192_reg_42434);

assign or_ln895_65_fu_36474_p2 = (xor_ln895_130_fu_36468_p2 | p_Result_195_reg_42465);

assign or_ln895_66_fu_36599_p2 = (xor_ln895_132_fu_36593_p2 | p_Result_198_reg_42496);

assign or_ln895_67_fu_36724_p2 = (xor_ln895_134_fu_36718_p2 | p_Result_201_reg_42527);

assign or_ln895_68_fu_33109_p2 = (xor_ln895_136_fu_33103_p2 | p_Result_204_fu_33025_p3);

assign or_ln895_69_fu_36866_p2 = (xor_ln895_138_fu_36860_p2 | p_Result_207_reg_42573);

assign or_ln895_6_fu_16957_p2 = (xor_ln895_12_fu_16951_p2 | p_Result_20_fu_16873_p3);

assign or_ln895_70_fu_36991_p2 = (xor_ln895_140_fu_36985_p2 | p_Result_210_reg_42604);

assign or_ln895_71_fu_37116_p2 = (xor_ln895_142_fu_37110_p2 | p_Result_213_reg_42635);

assign or_ln895_72_fu_37264_p2 = (xor_ln895_144_fu_37258_p2 | p_Result_216_fu_37193_p3);

assign or_ln895_73_fu_37413_p2 = (xor_ln895_146_fu_37407_p2 | p_Result_219_fu_37342_p3);

assign or_ln895_74_fu_37562_p2 = (xor_ln895_148_fu_37556_p2 | p_Result_222_fu_37491_p3);

assign or_ln895_75_fu_37711_p2 = (xor_ln895_150_fu_37705_p2 | p_Result_225_fu_37640_p3);

assign or_ln895_76_fu_33706_p2 = (xor_ln895_152_fu_33700_p2 | p_Result_228_fu_33622_p3);

assign or_ln895_77_fu_37877_p2 = (xor_ln895_154_fu_37871_p2 | p_Result_231_fu_37806_p3);

assign or_ln895_78_fu_38026_p2 = (xor_ln895_156_fu_38020_p2 | p_Result_234_fu_37955_p3);

assign or_ln895_79_fu_38175_p2 = (xor_ln895_158_fu_38169_p2 | p_Result_237_fu_38104_p3);

assign or_ln895_7_fu_19209_p2 = (xor_ln895_14_fu_19203_p2 | p_Result_23_reg_40525);

assign or_ln895_80_fu_38324_p2 = (xor_ln895_160_fu_38318_p2 | p_Result_240_fu_38253_p3);

assign or_ln895_8_fu_19333_p2 = (xor_ln895_16_fu_19327_p2 | p_Result_26_reg_40556);

assign or_ln895_9_fu_19481_p2 = (xor_ln895_18_fu_19475_p2 | p_Result_29_fu_19410_p3);

assign or_ln895_fu_18553_p2 = (xor_ln895_fu_18547_p2 | p_Result_2_reg_40340);

assign or_ln896_10_fu_17345_p2 = (xor_ln896_21_fu_17339_p2 | xor_ln896_20_fu_17245_p2);

assign or_ln896_11_fu_17489_p2 = (xor_ln896_23_fu_17483_p2 | xor_ln896_22_fu_17417_p2);

assign or_ln896_12_fu_19687_p2 = (xor_ln896_25_fu_19681_p2 | xor_ln896_24_fu_19601_p2);

assign or_ln896_13_fu_19836_p2 = (xor_ln896_27_fu_19830_p2 | xor_ln896_26_fu_19750_p2);

assign or_ln896_14_fu_17717_p2 = (xor_ln896_29_fu_17711_p2 | xor_ln896_28_fu_17645_p2);

assign or_ln896_15_fu_19978_p2 = (xor_ln896_31_fu_19972_p2 | xor_ln896_30_fu_19895_p2);

assign or_ln896_16_fu_20127_p2 = (xor_ln896_33_fu_20121_p2 | xor_ln896_32_fu_20041_p2);

assign or_ln896_17_fu_20276_p2 = (xor_ln896_35_fu_20270_p2 | xor_ln896_34_fu_20190_p2);

assign or_ln896_18_fu_20421_p2 = (xor_ln896_37_fu_20415_p2 | xor_ln896_36_fu_20335_p2);

assign or_ln896_19_fu_20550_p2 = (xor_ln896_39_fu_20544_p2 | xor_ln896_38_fu_20464_p2);

assign or_ln896_1_fu_18700_p2 = (xor_ln896_3_fu_18694_p2 | xor_ln896_2_fu_18617_p2);

assign or_ln896_20_fu_20683_p2 = (xor_ln896_41_fu_20677_p2 | xor_ln896_40_fu_20597_p2);

assign or_ln896_21_fu_20828_p2 = (xor_ln896_43_fu_20822_p2 | xor_ln896_42_fu_20742_p2);

assign or_ln896_22_fu_20957_p2 = (xor_ln896_45_fu_20951_p2 | xor_ln896_44_fu_20871_p2);

assign or_ln896_23_fu_21086_p2 = (xor_ln896_47_fu_21080_p2 | xor_ln896_46_fu_21000_p2);

assign or_ln896_24_fu_18355_p2 = (xor_ln896_49_fu_18349_p2 | xor_ln896_48_fu_18255_p2);

assign or_ln896_25_fu_21232_p2 = (xor_ln896_51_fu_21226_p2 | xor_ln896_50_fu_21146_p2);

assign or_ln896_26_fu_21361_p2 = (xor_ln896_53_fu_21355_p2 | xor_ln896_52_fu_21275_p2);

assign or_ln896_27_fu_24612_p2 = (xor_ln896_55_fu_24606_p2 | xor_ln896_54_fu_24529_p2);

assign or_ln896_28_fu_24736_p2 = (xor_ln896_57_fu_24730_p2 | xor_ln896_56_fu_24653_p2);

assign or_ln896_29_fu_24861_p2 = (xor_ln896_59_fu_24855_p2 | xor_ln896_58_fu_24778_p2);

assign or_ln896_2_fu_16603_p2 = (xor_ln896_5_fu_16597_p2 | xor_ln896_4_fu_16503_p2);

assign or_ln896_30_fu_24986_p2 = (xor_ln896_61_fu_24980_p2 | xor_ln896_60_fu_24903_p2);

assign or_ln896_31_fu_25111_p2 = (xor_ln896_63_fu_25105_p2 | xor_ln896_62_fu_25028_p2);

assign or_ln896_32_fu_25236_p2 = (xor_ln896_65_fu_25230_p2 | xor_ln896_64_fu_25153_p2);

assign or_ln896_33_fu_25361_p2 = (xor_ln896_67_fu_25355_p2 | xor_ln896_66_fu_25278_p2);

assign or_ln896_34_fu_25486_p2 = (xor_ln896_69_fu_25480_p2 | xor_ln896_68_fu_25403_p2);

assign or_ln896_35_fu_25608_p2 = (xor_ln896_71_fu_25602_p2 | xor_ln896_70_fu_25525_p2);

assign or_ln896_36_fu_25756_p2 = (xor_ln896_73_fu_25750_p2 | xor_ln896_72_fu_25670_p2);

assign or_ln896_37_fu_25905_p2 = (xor_ln896_75_fu_25899_p2 | xor_ln896_74_fu_25819_p2);

assign or_ln896_38_fu_26054_p2 = (xor_ln896_77_fu_26048_p2 | xor_ln896_76_fu_25968_p2);

assign or_ln896_39_fu_22304_p2 = (xor_ln896_79_fu_22298_p2 | xor_ln896_78_fu_22204_p2);

assign or_ln896_3_fu_18842_p2 = (xor_ln896_7_fu_18836_p2 | xor_ln896_6_fu_18759_p2);

assign or_ln896_40_fu_26220_p2 = (xor_ln896_81_fu_26214_p2 | xor_ln896_80_fu_26134_p2);

assign or_ln896_41_fu_26369_p2 = (xor_ln896_83_fu_26363_p2 | xor_ln896_82_fu_26283_p2);

assign or_ln896_42_fu_26518_p2 = (xor_ln896_85_fu_26512_p2 | xor_ln896_84_fu_26432_p2);

assign or_ln896_43_fu_26667_p2 = (xor_ln896_87_fu_26661_p2 | xor_ln896_86_fu_26581_p2);

assign or_ln896_44_fu_26816_p2 = (xor_ln896_89_fu_26810_p2 | xor_ln896_88_fu_26730_p2);

assign or_ln896_45_fu_27040_p2 = (xor_ln896_91_fu_27034_p2 | xor_ln896_90_fu_26940_p2);

assign or_ln896_46_fu_30716_p2 = (xor_ln896_93_fu_30710_p2 | xor_ln896_92_fu_30633_p2);

assign or_ln896_47_fu_30841_p2 = (xor_ln896_95_fu_30835_p2 | xor_ln896_94_fu_30758_p2);

assign or_ln896_48_fu_30966_p2 = (xor_ln896_97_fu_30960_p2 | xor_ln896_96_fu_30883_p2);

assign or_ln896_49_fu_31091_p2 = (xor_ln896_99_fu_31085_p2 | xor_ln896_98_fu_31008_p2);

assign or_ln896_4_fu_18967_p2 = (xor_ln896_9_fu_18961_p2 | xor_ln896_8_fu_18884_p2);

assign or_ln896_50_fu_31216_p2 = (xor_ln896_101_fu_31210_p2 | xor_ln896_100_fu_31133_p2);

assign or_ln896_51_fu_27574_p2 = (xor_ln896_103_fu_27568_p2 | xor_ln896_102_fu_27474_p2);

assign or_ln896_52_fu_31358_p2 = (xor_ln896_105_fu_31352_p2 | xor_ln896_104_fu_31275_p2);

assign or_ln896_53_fu_27835_p2 = (xor_ln896_107_fu_27829_p2 | xor_ln896_106_fu_27735_p2);

assign or_ln896_54_fu_31524_p2 = (xor_ln896_109_fu_31518_p2 | xor_ln896_108_fu_31438_p2);

assign or_ln896_55_fu_31673_p2 = (xor_ln896_111_fu_31667_p2 | xor_ln896_110_fu_31587_p2);

assign or_ln896_56_fu_31822_p2 = (xor_ln896_113_fu_31816_p2 | xor_ln896_112_fu_31736_p2);

assign or_ln896_57_fu_31971_p2 = (xor_ln896_115_fu_31965_p2 | xor_ln896_114_fu_31885_p2);

assign or_ln896_58_fu_32120_p2 = (xor_ln896_117_fu_32114_p2 | xor_ln896_116_fu_32034_p2);

assign or_ln896_59_fu_32269_p2 = (xor_ln896_119_fu_32263_p2 | xor_ln896_118_fu_32183_p2);

assign or_ln896_5_fu_19092_p2 = (xor_ln896_11_fu_19086_p2 | xor_ln896_10_fu_19009_p2);

assign or_ln896_60_fu_32418_p2 = (xor_ln896_121_fu_32412_p2 | xor_ln896_120_fu_32332_p2);

assign or_ln896_61_fu_28357_p2 = (xor_ln896_123_fu_28351_p2 | xor_ln896_122_fu_28257_p2);

assign or_ln896_62_fu_32584_p2 = (xor_ln896_125_fu_32578_p2 | xor_ln896_124_fu_32498_p2);

assign or_ln896_63_fu_36246_p2 = (xor_ln896_127_fu_36240_p2 | xor_ln896_126_fu_36163_p2);

assign or_ln896_64_fu_36371_p2 = (xor_ln896_129_fu_36365_p2 | xor_ln896_128_fu_36288_p2);

assign or_ln896_65_fu_36496_p2 = (xor_ln896_131_fu_36490_p2 | xor_ln896_130_fu_36413_p2);

assign or_ln896_66_fu_36621_p2 = (xor_ln896_133_fu_36615_p2 | xor_ln896_132_fu_36538_p2);

assign or_ln896_67_fu_36746_p2 = (xor_ln896_135_fu_36740_p2 | xor_ln896_134_fu_36663_p2);

assign or_ln896_68_fu_33133_p2 = (xor_ln896_137_fu_33127_p2 | xor_ln896_136_fu_33033_p2);

assign or_ln896_69_fu_36888_p2 = (xor_ln896_139_fu_36882_p2 | xor_ln896_138_fu_36805_p2);

assign or_ln896_6_fu_16981_p2 = (xor_ln896_13_fu_16975_p2 | xor_ln896_12_fu_16881_p2);

assign or_ln896_70_fu_37013_p2 = (xor_ln896_141_fu_37007_p2 | xor_ln896_140_fu_36930_p2);

assign or_ln896_71_fu_37138_p2 = (xor_ln896_143_fu_37132_p2 | xor_ln896_142_fu_37055_p2);

assign or_ln896_72_fu_37287_p2 = (xor_ln896_145_fu_37281_p2 | xor_ln896_144_fu_37201_p2);

assign or_ln896_73_fu_37436_p2 = (xor_ln896_147_fu_37430_p2 | xor_ln896_146_fu_37350_p2);

assign or_ln896_74_fu_37585_p2 = (xor_ln896_149_fu_37579_p2 | xor_ln896_148_fu_37499_p2);

assign or_ln896_75_fu_37734_p2 = (xor_ln896_151_fu_37728_p2 | xor_ln896_150_fu_37648_p2);

assign or_ln896_76_fu_33730_p2 = (xor_ln896_153_fu_33724_p2 | xor_ln896_152_fu_33630_p2);

assign or_ln896_77_fu_37900_p2 = (xor_ln896_155_fu_37894_p2 | xor_ln896_154_fu_37814_p2);

assign or_ln896_78_fu_38049_p2 = (xor_ln896_157_fu_38043_p2 | xor_ln896_156_fu_37963_p2);

assign or_ln896_79_fu_38198_p2 = (xor_ln896_159_fu_38192_p2 | xor_ln896_158_fu_38112_p2);

assign or_ln896_7_fu_19231_p2 = (xor_ln896_15_fu_19225_p2 | xor_ln896_14_fu_19148_p2);

assign or_ln896_80_fu_38347_p2 = (xor_ln896_161_fu_38341_p2 | xor_ln896_160_fu_38261_p2);

assign or_ln896_8_fu_19355_p2 = (xor_ln896_17_fu_19349_p2 | xor_ln896_16_fu_19272_p2);

assign or_ln896_9_fu_19504_p2 = (xor_ln896_19_fu_19498_p2 | xor_ln896_18_fu_19418_p2);

assign or_ln896_fu_18575_p2 = (xor_ln896_fu_18492_p2 | xor_ln896_1_fu_18569_p2);

assign overflow_100_fu_28563_p2 = (xor_ln895_181_fu_28557_p2 & p_Result_280_fu_28549_p3);

assign overflow_101_fu_28628_p2 = (xor_ln895_182_fu_28623_p2 & p_Result_282_reg_41729);

assign overflow_102_fu_28721_p2 = (xor_ln895_183_fu_28715_p2 & p_Result_284_fu_28707_p3);

assign overflow_103_fu_28821_p2 = (xor_ln895_184_fu_28815_p2 & p_Result_286_fu_28807_p3);

assign overflow_104_fu_28921_p2 = (xor_ln895_185_fu_28915_p2 & p_Result_288_fu_28907_p3);

assign overflow_105_fu_28986_p2 = (xor_ln895_186_fu_28981_p2 & p_Result_290_reg_41749);

assign overflow_106_fu_29079_p2 = (xor_ln895_187_fu_29073_p2 & p_Result_292_fu_29065_p3);

assign overflow_107_fu_29179_p2 = (xor_ln895_188_fu_29173_p2 & p_Result_294_fu_29165_p3);

assign overflow_108_fu_29281_p2 = (xor_ln895_189_fu_29275_p2 & p_Result_296_fu_29267_p3);

assign overflow_109_fu_29383_p2 = (xor_ln895_190_fu_29377_p2 & p_Result_298_fu_29369_p3);

assign overflow_10_fu_17333_p2 = (xor_ln895_21_fu_17327_p2 & or_ln895_10_fu_17321_p2);

assign overflow_110_fu_29485_p2 = (xor_ln895_191_fu_29479_p2 & p_Result_300_fu_29471_p3);

assign overflow_111_fu_29587_p2 = (xor_ln895_192_fu_29581_p2 & p_Result_302_fu_29573_p3);

assign overflow_112_fu_29689_p2 = (xor_ln895_193_fu_29683_p2 & p_Result_304_fu_29675_p3);

assign overflow_113_fu_29791_p2 = (xor_ln895_194_fu_29785_p2 & p_Result_306_fu_29777_p3);

assign overflow_114_fu_29893_p2 = (xor_ln895_195_fu_29887_p2 & p_Result_308_fu_29879_p3);

assign overflow_115_fu_29995_p2 = (xor_ln895_196_fu_29989_p2 & p_Result_310_fu_29981_p3);

assign overflow_116_fu_30097_p2 = (xor_ln895_197_fu_30091_p2 & p_Result_312_fu_30083_p3);

assign overflow_117_fu_33927_p2 = (xor_ln895_198_fu_33922_p2 & p_Result_314_reg_42247);

assign overflow_118_fu_33985_p2 = (xor_ln895_199_fu_33980_p2 & p_Result_316_reg_42267);

assign overflow_119_fu_30271_p2 = (xor_ln895_200_fu_30265_p2 & p_Result_318_fu_30257_p3);

assign overflow_11_fu_17477_p2 = (xor_ln895_21_fu_17327_p2 & or_ln895_11_fu_17471_p2);

assign overflow_120_fu_34043_p2 = (xor_ln895_201_fu_34038_p2 & p_Result_320_reg_42293);

assign overflow_121_fu_34101_p2 = (xor_ln895_202_fu_34096_p2 & p_Result_322_reg_42313);

assign overflow_122_fu_34159_p2 = (xor_ln895_203_fu_34154_p2 & p_Result_324_reg_42333);

assign overflow_123_fu_30481_p2 = (xor_ln895_204_fu_30475_p2 & p_Result_326_fu_30467_p3);

assign overflow_124_fu_34217_p2 = (xor_ln895_205_fu_34212_p2 & p_Result_328_reg_42359);

assign overflow_125_fu_34275_p2 = (xor_ln895_206_fu_34270_p2 & p_Result_330_reg_42379);

assign overflow_126_fu_34370_p2 = (xor_ln895_207_fu_34364_p2 & p_Result_332_fu_34356_p3);

assign overflow_127_fu_34472_p2 = (xor_ln895_208_fu_34466_p2 & p_Result_334_fu_34458_p3);

assign overflow_128_fu_34572_p2 = (xor_ln895_209_fu_34566_p2 & p_Result_336_fu_34558_p3);

assign overflow_129_fu_34674_p2 = (xor_ln895_210_fu_34668_p2 & p_Result_338_fu_34660_p3);

assign overflow_12_fu_19675_p2 = (xor_ln895_25_fu_19670_p2 & or_ln895_12_fu_19664_p2);

assign overflow_130_fu_34776_p2 = (xor_ln895_211_fu_34770_p2 & p_Result_340_fu_34762_p3);

assign overflow_131_fu_34878_p2 = (xor_ln895_212_fu_34872_p2 & p_Result_342_fu_34864_p3);

assign overflow_132_fu_34978_p2 = (xor_ln895_213_fu_34972_p2 & p_Result_344_fu_34964_p3);

assign overflow_133_fu_35080_p2 = (xor_ln895_214_fu_35074_p2 & p_Result_346_fu_35066_p3);

assign overflow_134_fu_35182_p2 = (xor_ln895_215_fu_35176_p2 & p_Result_348_fu_35168_p3);

assign overflow_135_fu_35284_p2 = (xor_ln895_216_fu_35278_p2 & p_Result_350_fu_35270_p3);

assign overflow_136_fu_35386_p2 = (xor_ln895_217_fu_35380_p2 & p_Result_352_fu_35372_p3);

assign overflow_137_fu_35488_p2 = (xor_ln895_218_fu_35482_p2 & p_Result_354_fu_35474_p3);

assign overflow_138_fu_35590_p2 = (xor_ln895_219_fu_35584_p2 & p_Result_356_fu_35576_p3);

assign overflow_139_fu_35692_p2 = (xor_ln895_220_fu_35686_p2 & p_Result_358_fu_35678_p3);

assign overflow_13_fu_19824_p2 = (xor_ln895_27_fu_19819_p2 & or_ln895_13_fu_19813_p2);

assign overflow_140_fu_35794_p2 = (xor_ln895_221_fu_35788_p2 & p_Result_360_fu_35780_p3);

assign overflow_141_fu_35896_p2 = (xor_ln895_222_fu_35890_p2 & p_Result_362_fu_35882_p3);

assign overflow_142_fu_35998_p2 = (xor_ln895_223_fu_35992_p2 & p_Result_364_fu_35984_p3);

assign overflow_143_fu_36100_p2 = (xor_ln895_224_fu_36094_p2 & p_Result_366_fu_36086_p3);

assign overflow_144_fu_38426_p2 = (xor_ln895_225_fu_38420_p2 & p_Result_368_fu_38412_p3);

assign overflow_145_fu_38526_p2 = (xor_ln895_226_fu_38520_p2 & p_Result_370_fu_38512_p3);

assign overflow_146_fu_38626_p2 = (xor_ln895_227_fu_38620_p2 & p_Result_372_fu_38612_p3);

assign overflow_147_fu_38726_p2 = (xor_ln895_228_fu_38720_p2 & p_Result_374_fu_38712_p3);

assign overflow_148_fu_38826_p2 = (xor_ln895_229_fu_38820_p2 & p_Result_376_fu_38812_p3);

assign overflow_149_fu_38926_p2 = (xor_ln895_230_fu_38920_p2 & p_Result_378_fu_38912_p3);

assign overflow_14_fu_17705_p2 = (xor_ln895_21_fu_17327_p2 & or_ln895_14_fu_17699_p2);

assign overflow_150_fu_39026_p2 = (xor_ln895_231_fu_39020_p2 & p_Result_380_fu_39012_p3);

assign overflow_151_fu_39126_p2 = (xor_ln895_232_fu_39120_p2 & p_Result_382_fu_39112_p3);

assign overflow_152_fu_39226_p2 = (xor_ln895_233_fu_39220_p2 & p_Result_384_fu_39212_p3);

assign overflow_153_fu_39328_p2 = (xor_ln895_234_fu_39322_p2 & p_Result_386_fu_39314_p3);

assign overflow_154_fu_39430_p2 = (xor_ln895_235_fu_39424_p2 & p_Result_388_fu_39416_p3);

assign overflow_155_fu_39532_p2 = (xor_ln895_236_fu_39526_p2 & p_Result_390_fu_39518_p3);

assign overflow_156_fu_39634_p2 = (xor_ln895_237_fu_39628_p2 & p_Result_392_fu_39620_p3);

assign overflow_157_fu_39736_p2 = (xor_ln895_238_fu_39730_p2 & p_Result_394_fu_39722_p3);

assign overflow_158_fu_39838_p2 = (xor_ln895_239_fu_39832_p2 & p_Result_396_fu_39824_p3);

assign overflow_159_fu_39940_p2 = (xor_ln895_240_fu_39934_p2 & p_Result_398_fu_39926_p3);

assign overflow_15_fu_19966_p2 = (xor_ln895_31_fu_19961_p2 & or_ln895_15_fu_19956_p2);

assign overflow_160_fu_40042_p2 = (xor_ln895_241_fu_40036_p2 & p_Result_400_fu_40028_p3);

assign overflow_161_fu_40144_p2 = (xor_ln895_242_fu_40138_p2 & p_Result_402_fu_40130_p3);

assign overflow_16_fu_20115_p2 = (xor_ln895_33_fu_20110_p2 & or_ln895_16_fu_20104_p2);

assign overflow_17_fu_20264_p2 = (xor_ln895_35_fu_20259_p2 & or_ln895_17_fu_20253_p2);

assign overflow_18_fu_20409_p2 = (xor_ln895_37_fu_20404_p2 & or_ln895_18_fu_20398_p2);

assign overflow_19_fu_20538_p2 = (xor_ln895_39_fu_20533_p2 & or_ln895_19_fu_20527_p2);

assign overflow_1_fu_18688_p2 = (xor_ln895_3_fu_18683_p2 & or_ln895_1_fu_18678_p2);

assign overflow_20_fu_20671_p2 = (xor_ln895_41_fu_20666_p2 & or_ln895_20_fu_20660_p2);

assign overflow_21_fu_20816_p2 = (xor_ln895_43_fu_20811_p2 & or_ln895_21_fu_20805_p2);

assign overflow_22_fu_20945_p2 = (xor_ln895_45_fu_20940_p2 & or_ln895_22_fu_20934_p2);

assign overflow_23_fu_21074_p2 = (xor_ln895_47_fu_21069_p2 & or_ln895_23_fu_21063_p2);

assign overflow_24_fu_18343_p2 = (xor_ln895_49_fu_18337_p2 & or_ln895_24_fu_18331_p2);

assign overflow_25_fu_21220_p2 = (xor_ln895_51_fu_21215_p2 & or_ln895_25_fu_21209_p2);

assign overflow_26_fu_21349_p2 = (xor_ln895_53_fu_21344_p2 & or_ln895_26_fu_21338_p2);

assign overflow_27_fu_24600_p2 = (xor_ln895_55_fu_24595_p2 & or_ln895_27_fu_24590_p2);

assign overflow_28_fu_24724_p2 = (xor_ln895_57_fu_24719_p2 & or_ln895_28_fu_24714_p2);

assign overflow_29_fu_24849_p2 = (xor_ln895_59_fu_24844_p2 & or_ln895_29_fu_24839_p2);

assign overflow_2_fu_16591_p2 = (xor_ln895_5_fu_16585_p2 & or_ln895_2_fu_16579_p2);

assign overflow_30_fu_24974_p2 = (xor_ln895_61_fu_24969_p2 & or_ln895_30_fu_24964_p2);

assign overflow_31_fu_25099_p2 = (xor_ln895_63_fu_25094_p2 & or_ln895_31_fu_25089_p2);

assign overflow_32_fu_25224_p2 = (xor_ln895_65_fu_25219_p2 & or_ln895_32_fu_25214_p2);

assign overflow_33_fu_25349_p2 = (xor_ln895_67_fu_25344_p2 & or_ln895_33_fu_25339_p2);

assign overflow_34_fu_25474_p2 = (xor_ln895_69_fu_25469_p2 & or_ln895_34_fu_25464_p2);

assign overflow_35_fu_25596_p2 = (xor_ln895_71_fu_25591_p2 & or_ln895_35_fu_25586_p2);

assign overflow_36_fu_25744_p2 = (xor_ln895_73_fu_25739_p2 & or_ln895_36_fu_25733_p2);

assign overflow_37_fu_25893_p2 = (xor_ln895_75_fu_25888_p2 & or_ln895_37_fu_25882_p2);

assign overflow_38_fu_26042_p2 = (xor_ln895_77_fu_26037_p2 & or_ln895_38_fu_26031_p2);

assign overflow_39_fu_22292_p2 = (xor_ln895_79_fu_22286_p2 & or_ln895_39_fu_22280_p2);

assign overflow_3_fu_18830_p2 = (xor_ln895_7_fu_18825_p2 & or_ln895_3_fu_18820_p2);

assign overflow_40_fu_26208_p2 = (xor_ln895_81_fu_26203_p2 & or_ln895_40_fu_26197_p2);

assign overflow_41_fu_26357_p2 = (xor_ln895_83_fu_26352_p2 & or_ln895_41_fu_26346_p2);

assign overflow_42_fu_26506_p2 = (xor_ln895_85_fu_26501_p2 & or_ln895_42_fu_26495_p2);

assign overflow_43_fu_26655_p2 = (xor_ln895_87_fu_26650_p2 & or_ln895_43_fu_26644_p2);

assign overflow_44_fu_26804_p2 = (xor_ln895_89_fu_26799_p2 & or_ln895_44_fu_26793_p2);

assign overflow_45_fu_27028_p2 = (xor_ln895_91_fu_27022_p2 & or_ln895_45_fu_27016_p2);

assign overflow_46_fu_30704_p2 = (xor_ln895_93_fu_30699_p2 & or_ln895_46_fu_30694_p2);

assign overflow_47_fu_30829_p2 = (xor_ln895_95_fu_30824_p2 & or_ln895_47_fu_30819_p2);

assign overflow_48_fu_30954_p2 = (xor_ln895_97_fu_30949_p2 & or_ln895_48_fu_30944_p2);

assign overflow_49_fu_31079_p2 = (xor_ln895_99_fu_31074_p2 & or_ln895_49_fu_31069_p2);

assign overflow_4_fu_18955_p2 = (xor_ln895_9_fu_18950_p2 & or_ln895_4_fu_18945_p2);

assign overflow_50_fu_31204_p2 = (xor_ln895_101_fu_31199_p2 & or_ln895_50_fu_31194_p2);

assign overflow_51_fu_27562_p2 = (xor_ln895_103_fu_27556_p2 & or_ln895_51_fu_27550_p2);

assign overflow_52_fu_31346_p2 = (xor_ln895_105_fu_31341_p2 & or_ln895_52_fu_31336_p2);

assign overflow_53_fu_27823_p2 = (xor_ln895_107_fu_27817_p2 & or_ln895_53_fu_27811_p2);

assign overflow_54_fu_31512_p2 = (xor_ln895_109_fu_31507_p2 & or_ln895_54_fu_31501_p2);

assign overflow_55_fu_31661_p2 = (xor_ln895_111_fu_31656_p2 & or_ln895_55_fu_31650_p2);

assign overflow_56_fu_31810_p2 = (xor_ln895_113_fu_31805_p2 & or_ln895_56_fu_31799_p2);

assign overflow_57_fu_31959_p2 = (xor_ln895_115_fu_31954_p2 & or_ln895_57_fu_31948_p2);

assign overflow_58_fu_32108_p2 = (xor_ln895_117_fu_32103_p2 & or_ln895_58_fu_32097_p2);

assign overflow_59_fu_32257_p2 = (xor_ln895_119_fu_32252_p2 & or_ln895_59_fu_32246_p2);

assign overflow_5_fu_19080_p2 = (xor_ln895_11_fu_19075_p2 & or_ln895_5_fu_19070_p2);

assign overflow_60_fu_32406_p2 = (xor_ln895_121_fu_32401_p2 & or_ln895_60_fu_32395_p2);

assign overflow_61_fu_28345_p2 = (xor_ln895_123_fu_28339_p2 & or_ln895_61_fu_28333_p2);

assign overflow_62_fu_32572_p2 = (xor_ln895_125_fu_32567_p2 & or_ln895_62_fu_32561_p2);

assign overflow_63_fu_36234_p2 = (xor_ln895_127_fu_36229_p2 & or_ln895_63_fu_36224_p2);

assign overflow_64_fu_36359_p2 = (xor_ln895_129_fu_36354_p2 & or_ln895_64_fu_36349_p2);

assign overflow_65_fu_36484_p2 = (xor_ln895_131_fu_36479_p2 & or_ln895_65_fu_36474_p2);

assign overflow_66_fu_36609_p2 = (xor_ln895_133_fu_36604_p2 & or_ln895_66_fu_36599_p2);

assign overflow_67_fu_36734_p2 = (xor_ln895_135_fu_36729_p2 & or_ln895_67_fu_36724_p2);

assign overflow_68_fu_33121_p2 = (xor_ln895_137_fu_33115_p2 & or_ln895_68_fu_33109_p2);

assign overflow_69_fu_36876_p2 = (xor_ln895_139_fu_36871_p2 & or_ln895_69_fu_36866_p2);

assign overflow_6_fu_16969_p2 = (xor_ln895_13_fu_16963_p2 & or_ln895_6_fu_16957_p2);

assign overflow_70_fu_37001_p2 = (xor_ln895_141_fu_36996_p2 & or_ln895_70_fu_36991_p2);

assign overflow_71_fu_37126_p2 = (xor_ln895_143_fu_37121_p2 & or_ln895_71_fu_37116_p2);

assign overflow_72_fu_37275_p2 = (xor_ln895_145_fu_37270_p2 & or_ln895_72_fu_37264_p2);

assign overflow_73_fu_37424_p2 = (xor_ln895_147_fu_37419_p2 & or_ln895_73_fu_37413_p2);

assign overflow_74_fu_37573_p2 = (xor_ln895_149_fu_37568_p2 & or_ln895_74_fu_37562_p2);

assign overflow_75_fu_37722_p2 = (xor_ln895_151_fu_37717_p2 & or_ln895_75_fu_37711_p2);

assign overflow_76_fu_33718_p2 = (xor_ln895_153_fu_33712_p2 & or_ln895_76_fu_33706_p2);

assign overflow_77_fu_37888_p2 = (xor_ln895_155_fu_37883_p2 & or_ln895_77_fu_37877_p2);

assign overflow_78_fu_38037_p2 = (xor_ln895_157_fu_38032_p2 & or_ln895_78_fu_38026_p2);

assign overflow_79_fu_38186_p2 = (xor_ln895_159_fu_38181_p2 & or_ln895_79_fu_38175_p2);

assign overflow_7_fu_19219_p2 = (xor_ln895_15_fu_19214_p2 & or_ln895_7_fu_19209_p2);

assign overflow_80_fu_38335_p2 = (xor_ln895_161_fu_38330_p2 & or_ln895_80_fu_38324_p2);

assign overflow_81_fu_22576_p2 = (xor_ln895_162_fu_22570_p2 & p_Result_242_fu_22562_p3);

assign overflow_82_fu_22674_p2 = (xor_ln895_163_fu_22668_p2 & p_Result_244_fu_22660_p3);

assign overflow_83_fu_22772_p2 = (xor_ln895_164_fu_22766_p2 & p_Result_246_fu_22758_p3);

assign overflow_84_fu_22870_p2 = (xor_ln895_165_fu_22864_p2 & p_Result_248_fu_22856_p3);

assign overflow_85_fu_22968_p2 = (xor_ln895_166_fu_22962_p2 & p_Result_250_fu_22954_p3);

assign overflow_86_fu_23066_p2 = (xor_ln895_167_fu_23060_p2 & p_Result_252_fu_23052_p3);

assign overflow_87_fu_23164_p2 = (xor_ln895_168_fu_23158_p2 & p_Result_254_fu_23150_p3);

assign overflow_88_fu_23262_p2 = (xor_ln895_169_fu_23256_p2 & p_Result_256_fu_23248_p3);

assign overflow_89_fu_23360_p2 = (xor_ln895_170_fu_23354_p2 & p_Result_258_fu_23346_p3);

assign overflow_8_fu_19343_p2 = (xor_ln895_17_fu_19338_p2 & or_ln895_8_fu_19333_p2);

assign overflow_90_fu_23462_p2 = (xor_ln895_171_fu_23456_p2 & p_Result_260_fu_23448_p3);

assign overflow_91_fu_23564_p2 = (xor_ln895_172_fu_23558_p2 & p_Result_262_fu_23550_p3);

assign overflow_92_fu_23666_p2 = (xor_ln895_173_fu_23660_p2 & p_Result_264_fu_23652_p3);

assign overflow_93_fu_23768_p2 = (xor_ln895_174_fu_23762_p2 & p_Result_266_fu_23754_p3);

assign overflow_94_fu_23870_p2 = (xor_ln895_175_fu_23864_p2 & p_Result_268_fu_23856_p3);

assign overflow_95_fu_23972_p2 = (xor_ln895_176_fu_23966_p2 & p_Result_270_fu_23958_p3);

assign overflow_96_fu_24074_p2 = (xor_ln895_177_fu_24068_p2 & p_Result_272_fu_24060_p3);

assign overflow_97_fu_24176_p2 = (xor_ln895_178_fu_24170_p2 & p_Result_274_fu_24162_p3);

assign overflow_98_fu_24278_p2 = (xor_ln895_179_fu_24272_p2 & p_Result_276_fu_24264_p3);

assign overflow_99_fu_28463_p2 = (xor_ln895_180_fu_28457_p2 & p_Result_278_fu_28449_p3);

assign overflow_9_fu_19492_p2 = (xor_ln895_19_fu_19487_p2 & or_ln895_9_fu_19481_p2);

assign overflow_fu_18563_p2 = (xor_ln895_1_fu_18558_p2 & or_ln895_fu_18553_p2);

assign p_Result_108_fu_25662_p3 = p_Val2_107_fu_25652_p2[32'd27];

assign p_Result_111_fu_25811_p3 = p_Val2_110_fu_25801_p2[32'd20];

assign p_Result_114_fu_25960_p3 = p_Val2_113_fu_25950_p2[32'd18];

assign p_Result_115_fu_22148_p3 = r_V_36_fu_22142_p2[32'd37];

assign p_Result_116_fu_22170_p3 = r_V_36_fu_22142_p2[32'd37];

assign p_Result_117_fu_22196_p3 = p_Val2_116_fu_22190_p2[32'd14];

assign p_Result_120_fu_26126_p3 = p_Val2_119_fu_26116_p2[32'd19];

assign p_Result_123_fu_26275_p3 = p_Val2_122_fu_26265_p2[32'd20];

assign p_Result_126_fu_26424_p3 = p_Val2_125_fu_26414_p2[32'd19];

assign p_Result_129_fu_26573_p3 = p_Val2_128_fu_26563_p2[32'd21];

assign p_Result_132_fu_26722_p3 = p_Val2_131_fu_26712_p2[32'd29];

assign p_Result_133_fu_26893_p3 = r_V_42_fu_26887_p2[32'd37];

assign p_Result_134_fu_26915_p3 = r_V_42_fu_26887_p2[32'd37];

assign p_Result_135_fu_26932_p3 = p_Val2_134_fu_26926_p2[32'd14];

assign p_Result_151_fu_27418_p3 = r_V_48_fu_27412_p2[32'd41];

assign p_Result_152_fu_27440_p3 = r_V_48_fu_27412_p2[32'd41];

assign p_Result_153_fu_27466_p3 = p_Val2_152_fu_27460_p2[32'd18];

assign p_Result_157_fu_27679_p3 = r_V_50_fu_27673_p2[32'd41];

assign p_Result_158_fu_27701_p3 = r_V_50_fu_27673_p2[32'd41];

assign p_Result_159_fu_27727_p3 = p_Val2_158_fu_27721_p2[32'd18];

assign p_Result_162_fu_31430_p3 = p_Val2_161_fu_31420_p2[32'd19];

assign p_Result_165_fu_31579_p3 = p_Val2_164_fu_31569_p2[32'd18];

assign p_Result_168_fu_31728_p3 = p_Val2_167_fu_31718_p2[32'd20];

assign p_Result_171_fu_31877_p3 = p_Val2_170_fu_31867_p2[32'd21];

assign p_Result_174_fu_32026_p3 = p_Val2_173_fu_32016_p2[32'd21];

assign p_Result_177_fu_32175_p3 = p_Val2_176_fu_32165_p2[32'd20];

assign p_Result_180_fu_32324_p3 = p_Val2_179_fu_32314_p2[32'd21];

assign p_Result_181_fu_28201_p3 = r_V_58_fu_28195_p2[32'd41];

assign p_Result_182_fu_28223_p3 = r_V_58_fu_28195_p2[32'd41];

assign p_Result_183_fu_28249_p3 = p_Val2_182_fu_28243_p2[32'd18];

assign p_Result_186_fu_32490_p3 = p_Val2_185_fu_32480_p2[32'd20];

assign p_Result_18_fu_16825_p3 = r_V_6_fu_16819_p2[32'd38];

assign p_Result_19_fu_16847_p3 = r_V_6_fu_16819_p2[32'd38];

assign p_Result_202_fu_32977_p3 = r_V_65_fu_32971_p2[32'd38];

assign p_Result_203_fu_32999_p3 = r_V_65_fu_32971_p2[32'd38];

assign p_Result_204_fu_33025_p3 = p_Val2_203_fu_33019_p2[32'd15];

assign p_Result_20_fu_16873_p3 = p_Val2_20_fu_16867_p2[32'd15];

assign p_Result_216_fu_37193_p3 = p_Val2_215_fu_37183_p2[32'd20];

assign p_Result_219_fu_37342_p3 = p_Val2_218_fu_37332_p2[32'd19];

assign p_Result_222_fu_37491_p3 = p_Val2_221_fu_37481_p2[32'd18];

assign p_Result_225_fu_37640_p3 = p_Val2_224_fu_37630_p2[32'd19];

assign p_Result_226_fu_33574_p3 = r_V_73_fu_33568_p2[32'd39];

assign p_Result_227_fu_33596_p3 = r_V_73_fu_33568_p2[32'd39];

assign p_Result_228_fu_33622_p3 = p_Val2_227_fu_33616_p2[32'd16];

assign p_Result_231_fu_37806_p3 = p_Val2_230_fu_37796_p2[32'd17];

assign p_Result_234_fu_37955_p3 = p_Val2_233_fu_37945_p2[32'd16];

assign p_Result_237_fu_38104_p3 = p_Val2_236_fu_38094_p2[32'd22];

assign p_Result_240_fu_38253_p3 = p_Val2_239_fu_38243_p2[32'd30];

assign p_Result_241_fu_22548_p3 = ret_V_fu_22542_p2[32'd32];

assign p_Result_242_fu_22562_p3 = p_Val2_241_fu_22556_p2[32'd31];

assign p_Result_243_fu_22646_p3 = ret_V_1_fu_22640_p2[32'd32];

assign p_Result_244_fu_22660_p3 = p_Val2_243_fu_22654_p2[32'd31];

assign p_Result_245_fu_22744_p3 = ret_V_2_fu_22738_p2[32'd32];

assign p_Result_246_fu_22758_p3 = p_Val2_245_fu_22752_p2[32'd31];

assign p_Result_247_fu_22842_p3 = ret_V_3_fu_22836_p2[32'd32];

assign p_Result_248_fu_22856_p3 = p_Val2_247_fu_22850_p2[32'd31];

assign p_Result_249_fu_22940_p3 = ret_V_4_fu_22934_p2[32'd32];

assign p_Result_250_fu_22954_p3 = p_Val2_249_fu_22948_p2[32'd31];

assign p_Result_251_fu_23038_p3 = ret_V_5_fu_23032_p2[32'd32];

assign p_Result_252_fu_23052_p3 = p_Val2_251_fu_23046_p2[32'd31];

assign p_Result_253_fu_23136_p3 = ret_V_6_fu_23130_p2[32'd32];

assign p_Result_254_fu_23150_p3 = p_Val2_253_fu_23144_p2[32'd31];

assign p_Result_255_fu_23234_p3 = ret_V_7_fu_23228_p2[32'd32];

assign p_Result_256_fu_23248_p3 = p_Val2_255_fu_23242_p2[32'd31];

assign p_Result_257_fu_23332_p3 = ret_V_8_fu_23326_p2[32'd32];

assign p_Result_258_fu_23346_p3 = p_Val2_257_fu_23340_p2[32'd31];

assign p_Result_259_fu_23434_p3 = ret_V_9_fu_23428_p2[32'd32];

assign p_Result_260_fu_23448_p3 = p_Val2_259_fu_23442_p2[32'd31];

assign p_Result_261_fu_23536_p3 = ret_V_10_fu_23530_p2[32'd32];

assign p_Result_262_fu_23550_p3 = p_Val2_261_fu_23544_p2[32'd31];

assign p_Result_263_fu_23638_p3 = ret_V_11_fu_23632_p2[32'd32];

assign p_Result_264_fu_23652_p3 = p_Val2_263_fu_23646_p2[32'd31];

assign p_Result_265_fu_23740_p3 = ret_V_12_fu_23734_p2[32'd32];

assign p_Result_266_fu_23754_p3 = p_Val2_265_fu_23748_p2[32'd31];

assign p_Result_267_fu_23842_p3 = ret_V_13_fu_23836_p2[32'd32];

assign p_Result_268_fu_23856_p3 = p_Val2_267_fu_23850_p2[32'd31];

assign p_Result_269_fu_23944_p3 = ret_V_14_fu_23938_p2[32'd32];

assign p_Result_270_fu_23958_p3 = p_Val2_269_fu_23952_p2[32'd31];

assign p_Result_271_fu_24046_p3 = ret_V_15_fu_24040_p2[32'd32];

assign p_Result_272_fu_24060_p3 = p_Val2_271_fu_24054_p2[32'd31];

assign p_Result_273_fu_24148_p3 = ret_V_16_fu_24142_p2[32'd32];

assign p_Result_274_fu_24162_p3 = p_Val2_273_fu_24156_p2[32'd31];

assign p_Result_275_fu_24250_p3 = ret_V_17_fu_24244_p2[32'd32];

assign p_Result_276_fu_24264_p3 = p_Val2_275_fu_24258_p2[32'd31];

assign p_Result_277_fu_28436_p3 = ret_V_18_fu_28430_p2[32'd32];

assign p_Result_278_fu_28449_p3 = p_Val2_277_fu_28444_p2[32'd31];

assign p_Result_279_fu_28536_p3 = ret_V_19_fu_28530_p2[32'd32];

assign p_Result_280_fu_28549_p3 = p_Val2_279_fu_28544_p2[32'd31];

assign p_Result_283_fu_28694_p3 = ret_V_21_fu_28688_p2[32'd32];

assign p_Result_284_fu_28707_p3 = p_Val2_283_fu_28702_p2[32'd31];

assign p_Result_285_fu_28794_p3 = ret_V_22_fu_28788_p2[32'd32];

assign p_Result_286_fu_28807_p3 = p_Val2_285_fu_28802_p2[32'd31];

assign p_Result_287_fu_28894_p3 = ret_V_23_fu_28888_p2[32'd32];

assign p_Result_288_fu_28907_p3 = p_Val2_287_fu_28902_p2[32'd31];

assign p_Result_291_fu_29052_p3 = ret_V_25_fu_29046_p2[32'd32];

assign p_Result_292_fu_29065_p3 = p_Val2_291_fu_29060_p2[32'd31];

assign p_Result_293_fu_29152_p3 = ret_V_26_fu_29146_p2[32'd32];

assign p_Result_294_fu_29165_p3 = p_Val2_293_fu_29160_p2[32'd31];

assign p_Result_295_fu_29253_p3 = ret_V_27_fu_29247_p2[32'd32];

assign p_Result_296_fu_29267_p3 = p_Val2_295_fu_29261_p2[32'd31];

assign p_Result_297_fu_29355_p3 = ret_V_28_fu_29349_p2[32'd32];

assign p_Result_298_fu_29369_p3 = p_Val2_297_fu_29363_p2[32'd31];

assign p_Result_299_fu_29457_p3 = ret_V_29_fu_29451_p2[32'd32];

assign p_Result_29_fu_19410_p3 = p_Val2_29_fu_19400_p2[32'd19];

assign p_Result_300_fu_29471_p3 = p_Val2_299_fu_29465_p2[32'd31];

assign p_Result_301_fu_29559_p3 = ret_V_30_fu_29553_p2[32'd32];

assign p_Result_302_fu_29573_p3 = p_Val2_301_fu_29567_p2[32'd31];

assign p_Result_303_fu_29661_p3 = ret_V_31_fu_29655_p2[32'd32];

assign p_Result_304_fu_29675_p3 = p_Val2_303_fu_29669_p2[32'd31];

assign p_Result_305_fu_29763_p3 = ret_V_32_fu_29757_p2[32'd32];

assign p_Result_306_fu_29777_p3 = p_Val2_305_fu_29771_p2[32'd31];

assign p_Result_307_fu_29865_p3 = ret_V_33_fu_29859_p2[32'd32];

assign p_Result_308_fu_29879_p3 = p_Val2_307_fu_29873_p2[32'd31];

assign p_Result_309_fu_29967_p3 = ret_V_34_fu_29961_p2[32'd32];

assign p_Result_30_fu_17189_p1 = p_read1_int_reg;

assign p_Result_30_fu_17189_p3 = p_Result_30_fu_17189_p1[32'd31];

assign p_Result_310_fu_29981_p3 = p_Val2_309_fu_29975_p2[32'd31];

assign p_Result_311_fu_30069_p3 = ret_V_35_fu_30063_p2[32'd32];

assign p_Result_312_fu_30083_p3 = p_Val2_311_fu_30077_p2[32'd31];

assign p_Result_317_fu_30243_p3 = ret_V_38_fu_30237_p2[32'd32];

assign p_Result_318_fu_30257_p3 = p_Val2_317_fu_30251_p2[32'd31];

assign p_Result_31_fu_17211_p1 = p_read1_int_reg;

assign p_Result_31_fu_17211_p3 = p_Result_31_fu_17211_p1[32'd31];

assign p_Result_325_fu_30453_p3 = ret_V_42_fu_30447_p2[32'd32];

assign p_Result_326_fu_30467_p3 = p_Val2_325_fu_30461_p2[32'd31];

assign p_Result_32_fu_17237_p3 = p_Val2_31_fu_17231_p2[32'd17];

assign p_Result_331_fu_34342_p3 = ret_V_45_fu_34336_p2[32'd32];

assign p_Result_332_fu_34356_p3 = p_Val2_331_fu_34350_p2[32'd31];

assign p_Result_333_fu_34444_p3 = ret_V_46_fu_34438_p2[32'd32];

assign p_Result_334_fu_34458_p3 = p_Val2_333_fu_34452_p2[32'd31];

assign p_Result_335_fu_34545_p3 = ret_V_47_fu_34539_p2[32'd32];

assign p_Result_336_fu_34558_p3 = p_Val2_335_fu_34553_p2[32'd31];

assign p_Result_337_fu_34646_p3 = ret_V_48_fu_34640_p2[32'd32];

assign p_Result_338_fu_34660_p3 = p_Val2_337_fu_34654_p2[32'd31];

assign p_Result_339_fu_34748_p3 = ret_V_49_fu_34742_p2[32'd32];

assign p_Result_33_fu_17383_p1 = p_read1_int_reg;

assign p_Result_33_fu_17383_p3 = p_Result_33_fu_17383_p1[32'd31];

assign p_Result_340_fu_34762_p3 = p_Val2_339_fu_34756_p2[32'd31];

assign p_Result_341_fu_34850_p3 = ret_V_50_fu_34844_p2[32'd32];

assign p_Result_342_fu_34864_p3 = p_Val2_341_fu_34858_p2[32'd31];

assign p_Result_343_fu_34951_p3 = ret_V_51_fu_34945_p2[32'd32];

assign p_Result_344_fu_34964_p3 = p_Val2_343_fu_34959_p2[32'd31];

assign p_Result_345_fu_35052_p3 = ret_V_52_fu_35046_p2[32'd32];

assign p_Result_346_fu_35066_p3 = p_Val2_345_fu_35060_p2[32'd31];

assign p_Result_347_fu_35154_p3 = ret_V_53_fu_35148_p2[32'd32];

assign p_Result_348_fu_35168_p3 = p_Val2_347_fu_35162_p2[32'd31];

assign p_Result_349_fu_35256_p3 = ret_V_54_fu_35250_p2[32'd32];

assign p_Result_34_fu_17409_p3 = p_Val2_33_fu_17403_p2[32'd13];

assign p_Result_350_fu_35270_p3 = p_Val2_349_fu_35264_p2[32'd31];

assign p_Result_351_fu_35358_p3 = ret_V_55_fu_35352_p2[32'd32];

assign p_Result_352_fu_35372_p3 = p_Val2_351_fu_35366_p2[32'd31];

assign p_Result_353_fu_35460_p3 = ret_V_56_fu_35454_p2[32'd32];

assign p_Result_354_fu_35474_p3 = p_Val2_353_fu_35468_p2[32'd31];

assign p_Result_355_fu_35562_p3 = ret_V_57_fu_35556_p2[32'd32];

assign p_Result_356_fu_35576_p3 = p_Val2_355_fu_35570_p2[32'd31];

assign p_Result_357_fu_35664_p3 = ret_V_58_fu_35658_p2[32'd32];

assign p_Result_358_fu_35678_p3 = p_Val2_357_fu_35672_p2[32'd31];

assign p_Result_359_fu_35766_p3 = ret_V_59_fu_35760_p2[32'd32];

assign p_Result_360_fu_35780_p3 = p_Val2_359_fu_35774_p2[32'd31];

assign p_Result_361_fu_35868_p3 = ret_V_60_fu_35862_p2[32'd32];

assign p_Result_362_fu_35882_p3 = p_Val2_361_fu_35876_p2[32'd31];

assign p_Result_363_fu_35970_p3 = ret_V_61_fu_35964_p2[32'd32];

assign p_Result_364_fu_35984_p3 = p_Val2_363_fu_35978_p2[32'd31];

assign p_Result_365_fu_36072_p3 = ret_V_62_fu_36066_p2[32'd32];

assign p_Result_366_fu_36086_p3 = p_Val2_365_fu_36080_p2[32'd31];

assign p_Result_367_fu_38399_p3 = ret_V_63_fu_38393_p2[32'd32];

assign p_Result_368_fu_38412_p3 = p_Val2_367_fu_38407_p2[32'd31];

assign p_Result_369_fu_38499_p3 = ret_V_64_fu_38493_p2[32'd32];

assign p_Result_370_fu_38512_p3 = p_Val2_369_fu_38507_p2[32'd31];

assign p_Result_371_fu_38599_p3 = ret_V_65_fu_38593_p2[32'd32];

assign p_Result_372_fu_38612_p3 = p_Val2_371_fu_38607_p2[32'd31];

assign p_Result_373_fu_38699_p3 = ret_V_66_fu_38693_p2[32'd32];

assign p_Result_374_fu_38712_p3 = p_Val2_373_fu_38707_p2[32'd31];

assign p_Result_375_fu_38799_p3 = ret_V_67_fu_38793_p2[32'd32];

assign p_Result_376_fu_38812_p3 = p_Val2_375_fu_38807_p2[32'd31];

assign p_Result_377_fu_38899_p3 = ret_V_68_fu_38893_p2[32'd32];

assign p_Result_378_fu_38912_p3 = p_Val2_377_fu_38907_p2[32'd31];

assign p_Result_379_fu_38999_p3 = ret_V_69_fu_38993_p2[32'd32];

assign p_Result_37_fu_19593_p3 = p_Val2_36_fu_19583_p2[32'd21];

assign p_Result_380_fu_39012_p3 = p_Val2_379_fu_39007_p2[32'd31];

assign p_Result_381_fu_39099_p3 = ret_V_70_fu_39093_p2[32'd32];

assign p_Result_382_fu_39112_p3 = p_Val2_381_fu_39107_p2[32'd31];

assign p_Result_383_fu_39199_p3 = ret_V_71_fu_39193_p2[32'd32];

assign p_Result_384_fu_39212_p3 = p_Val2_383_fu_39207_p2[32'd31];

assign p_Result_385_fu_39300_p3 = ret_V_72_fu_39294_p2[32'd32];

assign p_Result_386_fu_39314_p3 = p_Val2_385_fu_39308_p2[32'd31];

assign p_Result_387_fu_39402_p3 = ret_V_73_fu_39396_p2[32'd32];

assign p_Result_388_fu_39416_p3 = p_Val2_387_fu_39410_p2[32'd31];

assign p_Result_389_fu_39504_p3 = ret_V_74_fu_39498_p2[32'd32];

assign p_Result_390_fu_39518_p3 = p_Val2_389_fu_39512_p2[32'd31];

assign p_Result_391_fu_39606_p3 = ret_V_75_fu_39600_p2[32'd32];

assign p_Result_392_fu_39620_p3 = p_Val2_391_fu_39614_p2[32'd31];

assign p_Result_393_fu_39708_p3 = ret_V_76_fu_39702_p2[32'd32];

assign p_Result_394_fu_39722_p3 = p_Val2_393_fu_39716_p2[32'd31];

assign p_Result_395_fu_39810_p3 = ret_V_77_fu_39804_p2[32'd32];

assign p_Result_396_fu_39824_p3 = p_Val2_395_fu_39818_p2[32'd31];

assign p_Result_397_fu_39912_p3 = ret_V_78_fu_39906_p2[32'd32];

assign p_Result_398_fu_39926_p3 = p_Val2_397_fu_39920_p2[32'd31];

assign p_Result_399_fu_40014_p3 = ret_V_79_fu_40008_p2[32'd32];

assign p_Result_400_fu_40028_p3 = p_Val2_399_fu_40022_p2[32'd31];

assign p_Result_401_fu_40116_p3 = ret_V_80_fu_40110_p2[32'd32];

assign p_Result_402_fu_40130_p3 = p_Val2_401_fu_40124_p2[32'd31];

assign p_Result_40_fu_19742_p3 = p_Val2_39_fu_19732_p2[32'd21];

assign p_Result_41_fu_17611_p1 = p_read1_int_reg;

assign p_Result_41_fu_17611_p3 = p_Result_41_fu_17611_p1[32'd31];

assign p_Result_42_fu_17637_p3 = p_Val2_41_fu_17631_p2[32'd16];

assign p_Result_48_fu_20033_p3 = p_Val2_47_fu_20023_p2[32'd19];

assign p_Result_51_fu_20182_p3 = p_Val2_50_fu_20172_p2[32'd21];

assign p_Result_54_fu_20327_p3 = p_Val2_53_fu_20321_p2[32'd19];

assign p_Result_57_fu_20456_p3 = p_Val2_56_fu_20450_p2[32'd20];

assign p_Result_60_fu_20589_p3 = p_Val2_59_fu_20579_p2[32'd18];

assign p_Result_63_fu_20734_p3 = p_Val2_62_fu_20728_p2[32'd19];

assign p_Result_66_fu_20863_p3 = p_Val2_65_fu_20857_p2[32'd19];

assign p_Result_69_fu_20992_p3 = p_Val2_68_fu_20986_p2[32'd14];

assign p_Result_6_fu_16441_p3 = r_V_2_fu_16435_p2[32'd38];

assign p_Result_70_fu_18199_p3 = r_V_21_fu_18193_p2[32'd38];

assign p_Result_71_fu_18221_p3 = r_V_21_fu_18193_p2[32'd38];

assign p_Result_72_fu_18247_p3 = p_Val2_71_fu_18241_p2[32'd15];

assign p_Result_75_fu_21138_p3 = p_Val2_74_fu_21132_p2[32'd21];

assign p_Result_78_fu_21267_p3 = p_Val2_77_fu_21261_p2[32'd19];

assign p_Result_7_fu_16469_p3 = r_V_2_fu_16435_p2[32'd38];

assign p_Result_8_fu_16495_p3 = p_Val2_8_fu_16489_p2[32'd15];

assign p_Val2_100_fu_21860_p4 = {{r_V_31_fu_496_p2[45:24]}};

assign p_Val2_101_fu_21894_p2 = ($signed(zext_ln377_34_fu_21890_p1) + $signed(sext_ln823_32_fu_21870_p1));

assign p_Val2_103_fu_21924_p4 = {{r_V_32_fu_499_p2[55:24]}};

assign p_Val2_104_fu_21954_p2 = (zext_ln377_35_fu_21950_p1 + p_Val2_103_fu_21924_p4);

assign p_Val2_107_fu_25652_p2 = ($signed(zext_ln377_36_fu_25649_p1) + $signed(sext_ln823_33_fu_25646_p1));

assign p_Val2_10_fu_16635_p4 = {{r_V_3_fu_510_p2[44:24]}};

assign p_Val2_110_fu_25801_p2 = ($signed(zext_ln377_37_fu_25798_p1) + $signed(sext_ln823_34_fu_25795_p1));

assign p_Val2_113_fu_25950_p2 = ($signed(zext_ln377_38_fu_25947_p1) + $signed(sext_ln823_35_fu_25944_p1));

assign p_Val2_115_fu_22156_p4 = {{r_V_36_fu_22142_p2[37:24]}};

assign p_Val2_116_fu_22190_p2 = ($signed(zext_ln377_39_fu_22186_p1) + $signed(sext_ln823_36_fu_22166_p1));

assign p_Val2_119_fu_26116_p2 = ($signed(zext_ln377_40_fu_26113_p1) + $signed(sext_ln823_37_fu_26110_p1));

assign p_Val2_11_fu_16669_p2 = ($signed(zext_ln377_3_fu_16665_p1) + $signed(sext_ln823_6_fu_16645_p1));

assign p_Val2_122_fu_26265_p2 = ($signed(zext_ln377_41_fu_26262_p1) + $signed(sext_ln823_38_fu_26259_p1));

assign p_Val2_125_fu_26414_p2 = ($signed(zext_ln377_42_fu_26411_p1) + $signed(sext_ln823_39_fu_26408_p1));

assign p_Val2_128_fu_26563_p2 = ($signed(zext_ln377_43_fu_26560_p1) + $signed(sext_ln823_40_fu_26557_p1));

assign p_Val2_131_fu_26712_p2 = ($signed(zext_ln377_44_fu_26709_p1) + $signed(sext_ln823_41_fu_26706_p1));

assign p_Val2_133_fu_26901_p4 = {{r_V_42_fu_26887_p2[37:24]}};

assign p_Val2_134_fu_26926_p2 = ($signed(zext_ln377_45_fu_26923_p1) + $signed(sext_ln823_42_fu_26911_p1));

assign p_Val2_136_fu_27072_p4 = {{r_V_43_fu_531_p2[42:24]}};

assign p_Val2_137_fu_27106_p2 = ($signed(zext_ln377_46_fu_27102_p1) + $signed(sext_ln823_43_fu_27082_p1));

assign p_Val2_139_fu_27136_p4 = {{r_V_44_fu_520_p2[41:24]}};

assign p_Val2_13_fu_16699_p4 = {{r_V_4_fu_526_p2[42:24]}};

assign p_Val2_140_fu_27170_p2 = ($signed(zext_ln377_47_fu_27166_p1) + $signed(sext_ln823_44_fu_27146_p1));

assign p_Val2_142_fu_27200_p4 = {{r_V_45_fu_506_p2[44:24]}};

assign p_Val2_143_fu_27234_p2 = ($signed(zext_ln377_48_fu_27230_p1) + $signed(sext_ln823_45_fu_27210_p1));

assign p_Val2_145_fu_27264_p4 = {{r_V_46_fu_530_p2[43:24]}};

assign p_Val2_146_fu_27298_p2 = ($signed(zext_ln377_49_fu_27294_p1) + $signed(sext_ln823_46_fu_27274_p1));

assign p_Val2_148_fu_27328_p4 = {{r_V_47_fu_471_p2[42:24]}};

assign p_Val2_149_fu_27362_p2 = ($signed(zext_ln377_50_fu_27358_p1) + $signed(sext_ln823_47_fu_27338_p1));

assign p_Val2_14_fu_16733_p2 = ($signed(zext_ln377_4_fu_16729_p1) + $signed(sext_ln823_7_fu_16709_p1));

assign p_Val2_151_fu_27426_p4 = {{r_V_48_fu_27412_p2[41:24]}};

assign p_Val2_152_fu_27460_p2 = ($signed(zext_ln377_51_fu_27456_p1) + $signed(sext_ln823_48_fu_27436_p1));

assign p_Val2_154_fu_27606_p4 = {{r_V_49_fu_480_p2[42:24]}};

assign p_Val2_155_fu_27640_p2 = ($signed(zext_ln377_52_fu_27636_p1) + $signed(sext_ln823_49_fu_27616_p1));

assign p_Val2_157_fu_27687_p4 = {{r_V_50_fu_27673_p2[41:24]}};

assign p_Val2_158_fu_27721_p2 = ($signed(zext_ln377_53_fu_27717_p1) + $signed(sext_ln823_50_fu_27697_p1));

assign p_Val2_161_fu_31420_p2 = ($signed(zext_ln377_54_fu_31417_p1) + $signed(sext_ln823_51_fu_31414_p1));

assign p_Val2_164_fu_31569_p2 = ($signed(zext_ln377_55_fu_31566_p1) + $signed(sext_ln823_52_fu_31563_p1));

assign p_Val2_167_fu_31718_p2 = ($signed(zext_ln377_56_fu_31715_p1) + $signed(sext_ln823_53_fu_31712_p1));

assign p_Val2_16_fu_16763_p4 = {{r_V_5_fu_500_p2[42:24]}};

assign p_Val2_170_fu_31867_p2 = ($signed(zext_ln377_57_fu_31864_p1) + $signed(sext_ln823_54_fu_31861_p1));

assign p_Val2_173_fu_32016_p2 = ($signed(zext_ln377_58_fu_32013_p1) + $signed(sext_ln823_55_fu_32010_p1));

assign p_Val2_176_fu_32165_p2 = ($signed(zext_ln377_59_fu_32162_p1) + $signed(sext_ln823_56_fu_32159_p1));

assign p_Val2_179_fu_32314_p2 = ($signed(zext_ln377_60_fu_32311_p1) + $signed(sext_ln823_57_fu_32308_p1));

assign p_Val2_17_fu_16797_p2 = ($signed(zext_ln377_5_fu_16793_p1) + $signed(sext_ln823_8_fu_16773_p1));

assign p_Val2_181_fu_28209_p4 = {{r_V_58_fu_28195_p2[41:24]}};

assign p_Val2_182_fu_28243_p2 = ($signed(zext_ln377_61_fu_28239_p1) + $signed(sext_ln823_58_fu_28219_p1));

assign p_Val2_185_fu_32480_p2 = ($signed(zext_ln377_62_fu_32477_p1) + $signed(sext_ln823_59_fu_32474_p1));

assign p_Val2_187_fu_32648_p4 = {{r_V_60_fu_474_p2[41:24]}};

assign p_Val2_188_fu_32682_p2 = ($signed(zext_ln377_63_fu_32678_p1) + $signed(sext_ln823_60_fu_32658_p1));

assign p_Val2_190_fu_32712_p4 = {{r_V_61_fu_543_p2[42:24]}};

assign p_Val2_191_fu_32746_p2 = ($signed(zext_ln377_64_fu_32742_p1) + $signed(sext_ln823_61_fu_32722_p1));

assign p_Val2_193_fu_32776_p4 = {{r_V_62_fu_477_p2[43:24]}};

assign p_Val2_194_fu_32810_p2 = ($signed(zext_ln377_65_fu_32806_p1) + $signed(sext_ln823_62_fu_32786_p1));

assign p_Val2_196_fu_32840_p4 = {{r_V_63_fu_545_p2[41:24]}};

assign p_Val2_197_fu_32874_p2 = ($signed(zext_ln377_66_fu_32870_p1) + $signed(sext_ln823_63_fu_32850_p1));

assign p_Val2_199_fu_32904_p4 = {{r_V_64_fu_533_p2[43:24]}};

assign p_Val2_19_fu_16833_p4 = {{r_V_6_fu_16819_p2[38:24]}};

assign p_Val2_1_fu_16291_p4 = {{r_V_fu_519_p2[46:24]}};

assign p_Val2_200_fu_32938_p2 = ($signed(zext_ln377_67_fu_32934_p1) + $signed(sext_ln823_64_fu_32914_p1));

assign p_Val2_202_fu_32985_p4 = {{r_V_65_fu_32971_p2[38:24]}};

assign p_Val2_203_fu_33019_p2 = ($signed(zext_ln377_68_fu_33015_p1) + $signed(sext_ln823_65_fu_32995_p1));

assign p_Val2_205_fu_33165_p4 = {{r_V_66_fu_511_p2[42:24]}};

assign p_Val2_206_fu_33199_p2 = ($signed(zext_ln377_69_fu_33195_p1) + $signed(sext_ln823_66_fu_33175_p1));

assign p_Val2_208_fu_33229_p4 = {{r_V_67_fu_522_p2[43:24]}};

assign p_Val2_209_fu_33263_p2 = ($signed(zext_ln377_70_fu_33259_p1) + $signed(sext_ln823_67_fu_33239_p1));

assign p_Val2_20_fu_16867_p2 = ($signed(zext_ln377_6_fu_16863_p1) + $signed(sext_ln823_9_fu_16843_p1));

assign p_Val2_211_fu_33293_p4 = {{r_V_68_fu_544_p2[41:24]}};

assign p_Val2_212_fu_33327_p2 = ($signed(zext_ln377_71_fu_33323_p1) + $signed(sext_ln823_68_fu_33303_p1));

assign p_Val2_215_fu_37183_p2 = ($signed(zext_ln377_72_fu_37180_p1) + $signed(sext_ln823_69_fu_37177_p1));

assign p_Val2_218_fu_37332_p2 = ($signed(zext_ln377_73_fu_37329_p1) + $signed(sext_ln823_70_fu_37326_p1));

assign p_Val2_221_fu_37481_p2 = ($signed(zext_ln377_74_fu_37478_p1) + $signed(sext_ln823_71_fu_37475_p1));

assign p_Val2_224_fu_37630_p2 = ($signed(zext_ln377_75_fu_37627_p1) + $signed(sext_ln823_72_fu_37624_p1));

assign p_Val2_226_fu_33582_p4 = {{r_V_73_fu_33568_p2[39:24]}};

assign p_Val2_227_fu_33616_p2 = ($signed(zext_ln377_76_fu_33612_p1) + $signed(sext_ln823_73_fu_33592_p1));

assign p_Val2_22_fu_17013_p4 = {{r_V_7_fu_537_p2[55:24]}};

assign p_Val2_230_fu_37796_p2 = ($signed(zext_ln377_77_fu_37793_p1) + $signed(sext_ln823_74_fu_37790_p1));

assign p_Val2_233_fu_37945_p2 = ($signed(zext_ln377_78_fu_37942_p1) + $signed(sext_ln823_75_fu_37939_p1));

assign p_Val2_236_fu_38094_p2 = ($signed(zext_ln377_79_fu_38091_p1) + $signed(sext_ln823_76_fu_38088_p1));

assign p_Val2_239_fu_38243_p2 = ($signed(zext_ln377_80_fu_38240_p1) + $signed(sext_ln823_77_fu_38237_p1));

assign p_Val2_23_fu_17043_p2 = (zext_ln377_7_fu_17039_p1 + p_Val2_22_fu_17013_p4);

assign p_Val2_241_fu_22556_p2 = ($signed(rhs_fu_18606_p3) + $signed(32'd140968));

assign p_Val2_243_fu_22654_p2 = ($signed(rhs_1_fu_18731_p3) + $signed(32'd4294771000));

assign p_Val2_245_fu_22752_p2 = ($signed(rhs_2_fu_18749_p3) + $signed(32'd4293355132));

assign p_Val2_247_fu_22850_p2 = ($signed(rhs_3_fu_18873_p3) + $signed(32'd4293905382));

assign p_Val2_249_fu_22948_p2 = ($signed(rhs_4_fu_18998_p3) + $signed(32'd4294962961));

assign p_Val2_251_fu_23046_p2 = ($signed(rhs_5_fu_19123_p3) + $signed(32'd4294961617));

assign p_Val2_253_fu_23144_p2 = ($signed(rhs_6_fu_19141_p3) + $signed(32'd4294940721));

assign p_Val2_255_fu_23242_p2 = ($signed(rhs_7_fu_19262_p3) + $signed(32'd5062185));

assign p_Val2_257_fu_23340_p2 = ($signed(rhs_8_fu_19386_p3) + $signed(32'd6923874));

assign p_Val2_259_fu_23442_p2 = ($signed(rhs_9_fu_19535_p3) + $signed(lhs_fu_22628_p3));

assign p_Val2_25_fu_17073_p4 = {{r_V_8_fu_514_p2[44:24]}};

assign p_Val2_261_fu_23544_p2 = ($signed(rhs_10_fu_19553_p3) + $signed(lhs_1_fu_22726_p3));

assign p_Val2_263_fu_23646_p2 = ($signed(rhs_11_fu_19570_p3) + $signed(lhs_2_fu_22824_p3));

assign p_Val2_265_fu_23748_p2 = ($signed(rhs_12_fu_19718_p3) + $signed(lhs_3_fu_22922_p3));

assign p_Val2_267_fu_23850_p2 = ($signed(rhs_13_fu_19867_p3) + $signed(lhs_4_fu_23020_p3));

assign p_Val2_269_fu_23952_p2 = ($signed(rhs_14_fu_19885_p3) + $signed(lhs_5_fu_23118_p3));

assign p_Val2_26_fu_17107_p2 = ($signed(zext_ln377_8_fu_17103_p1) + $signed(sext_ln823_10_fu_17083_p1));

assign p_Val2_271_fu_24054_p2 = ($signed(rhs_15_fu_20009_p3) + $signed(lhs_6_fu_23216_p3));

assign p_Val2_273_fu_24156_p2 = ($signed(rhs_16_fu_20158_p3) + $signed(lhs_7_fu_23314_p3));

assign p_Val2_275_fu_24258_p2 = ($signed(rhs_17_fu_20307_p3) + $signed(lhs_8_fu_23412_p3));

assign p_Val2_277_fu_28444_p2 = ($signed(rhs_18_fu_24420_p3) + $signed(lhs_9_reg_41674));

assign p_Val2_279_fu_28544_p2 = ($signed(rhs_19_fu_24437_p3) + $signed(lhs_10_reg_41680));

assign p_Val2_281_fu_24360_p2 = ($signed(rhs_20_fu_20714_p3) + $signed(lhs_11_fu_23718_p3));

assign p_Val2_283_fu_28702_p2 = ($signed(rhs_21_fu_24454_p3) + $signed(lhs_12_reg_41686));

assign p_Val2_285_fu_28802_p2 = ($signed(rhs_22_fu_24471_p3) + $signed(lhs_13_reg_41692));

assign p_Val2_287_fu_28902_p2 = ($signed(rhs_23_fu_24488_p3) + $signed(lhs_14_reg_41698));

assign p_Val2_289_fu_24396_p2 = ($signed(rhs_24_fu_21119_p3) + $signed(lhs_15_fu_24126_p3));

assign p_Val2_291_fu_29060_p2 = ($signed(rhs_25_fu_24505_p3) + $signed(lhs_16_reg_41704));

assign p_Val2_293_fu_29160_p2 = ($signed(rhs_26_fu_24522_p3) + $signed(lhs_17_reg_41710));

assign p_Val2_295_fu_29261_p2 = ($signed(rhs_27_fu_24643_p3) + $signed(lhs_18_fu_28515_p3));

assign p_Val2_297_fu_29363_p2 = ($signed(rhs_28_fu_24767_p3) + $signed(lhs_19_fu_28615_p3));

assign p_Val2_299_fu_29465_p2 = ($signed(rhs_29_fu_24892_p3) + $signed(lhs_20_fu_28673_p3));

assign p_Val2_29_fu_19400_p2 = ($signed(zext_ln377_9_fu_19397_p1) + $signed(sext_ln823_11_fu_19394_p1));

assign p_Val2_2_fu_16325_p2 = ($signed(zext_ln377_fu_16321_p1) + $signed(sext_ln823_3_fu_16301_p1));

assign p_Val2_301_fu_29567_p2 = ($signed(rhs_30_fu_25017_p3) + $signed(lhs_21_fu_28773_p3));

assign p_Val2_303_fu_29669_p2 = ($signed(rhs_31_fu_25142_p3) + $signed(lhs_22_fu_28873_p3));

assign p_Val2_305_fu_29771_p2 = ($signed(rhs_32_fu_25267_p3) + $signed(lhs_23_fu_28973_p3));

assign p_Val2_307_fu_29873_p2 = ($signed(rhs_33_fu_25392_p3) + $signed(lhs_24_fu_29031_p3));

assign p_Val2_309_fu_29975_p2 = ($signed(rhs_34_fu_25517_p3) + $signed(lhs_25_fu_29131_p3));

assign p_Val2_30_fu_17197_p1 = p_read1_int_reg;

assign p_Val2_30_fu_17197_p4 = {{p_Val2_30_fu_17197_p1[31:15]}};

assign p_Val2_311_fu_30077_p2 = ($signed(rhs_35_fu_25639_p3) + $signed(lhs_26_fu_29231_p3));

assign p_Val2_313_fu_30179_p2 = ($signed(rhs_36_fu_25787_p3) + $signed(lhs_27_fu_29333_p3));

assign p_Val2_315_fu_30215_p2 = ($signed(rhs_37_fu_25936_p3) + $signed(lhs_28_fu_29435_p3));

assign p_Val2_317_fu_30251_p2 = ($signed(rhs_38_fu_26085_p3) + $signed(lhs_29_fu_29537_p3));

assign p_Val2_319_fu_30353_p2 = ($signed(rhs_39_fu_26103_p3) + $signed(lhs_30_fu_29639_p3));

assign p_Val2_31_fu_17231_p2 = ($signed(zext_ln377_10_fu_17227_p1) + $signed(sext_ln823_fu_17207_p1));

assign p_Val2_321_fu_30389_p2 = ($signed(rhs_40_fu_26251_p3) + $signed(lhs_31_fu_29741_p3));

assign p_Val2_323_fu_30425_p2 = ($signed(rhs_41_fu_26400_p3) + $signed(lhs_32_fu_29843_p3));

assign p_Val2_325_fu_30461_p2 = ($signed(rhs_42_fu_26549_p3) + $signed(lhs_33_fu_29945_p3));

assign p_Val2_327_fu_30563_p2 = ($signed(rhs_43_fu_26698_p3) + $signed(lhs_34_fu_30047_p3));

assign p_Val2_329_fu_30599_p2 = ($signed(rhs_44_fu_26847_p3) + $signed(lhs_35_fu_30149_p3));

assign p_Val2_32_fu_17369_p1 = p_read1_int_reg;

assign p_Val2_32_fu_17369_p4 = {{p_Val2_32_fu_17369_p1[31:19]}};

assign p_Val2_331_fu_34350_p2 = ($signed(rhs_45_fu_30623_p3) + $signed(lhs_36_fu_33972_p3));

assign p_Val2_333_fu_34452_p2 = ($signed(rhs_46_fu_30747_p3) + $signed(lhs_37_fu_34030_p3));

assign p_Val2_335_fu_34553_p2 = ($signed(rhs_47_fu_30872_p3) + $signed(lhs_38_reg_42274));

assign p_Val2_337_fu_34654_p2 = ($signed(rhs_48_fu_30997_p3) + $signed(lhs_39_fu_34088_p3));

assign p_Val2_339_fu_34756_p2 = ($signed(rhs_49_fu_31122_p3) + $signed(lhs_40_fu_34146_p3));

assign p_Val2_33_fu_17403_p2 = ($signed(zext_ln377_11_fu_17399_p1) + $signed(sext_ln823_1_fu_17379_p1));

assign p_Val2_341_fu_34858_p2 = ($signed(rhs_50_fu_31247_p3) + $signed(lhs_41_fu_34204_p3));

assign p_Val2_343_fu_34959_p2 = ($signed(rhs_51_fu_31265_p3) + $signed(lhs_42_reg_42340));

assign p_Val2_345_fu_35060_p2 = ($signed(rhs_52_fu_31389_p3) + $signed(lhs_43_fu_34262_p3));

assign p_Val2_347_fu_35162_p2 = ($signed(rhs_53_fu_31407_p3) + $signed(lhs_44_fu_34320_p3));

assign p_Val2_349_fu_35264_p2 = ($signed(rhs_54_fu_31555_p3) + $signed(lhs_45_fu_34422_p3));

assign p_Val2_351_fu_35366_p2 = ($signed(rhs_55_fu_31704_p3) + $signed(lhs_46_fu_34524_p3));

assign p_Val2_353_fu_35468_p2 = ($signed(rhs_56_fu_31853_p3) + $signed(lhs_47_fu_34624_p3));

assign p_Val2_355_fu_35570_p2 = ($signed(rhs_57_fu_32002_p3) + $signed(lhs_48_fu_34726_p3));

assign p_Val2_357_fu_35672_p2 = ($signed(rhs_58_fu_32151_p3) + $signed(lhs_49_fu_34828_p3));

assign p_Val2_359_fu_35774_p2 = ($signed(rhs_59_fu_32300_p3) + $signed(lhs_50_fu_34930_p3));

assign p_Val2_361_fu_35876_p2 = ($signed(rhs_60_fu_32449_p3) + $signed(lhs_51_fu_35030_p3));

assign p_Val2_363_fu_35978_p2 = ($signed(rhs_61_fu_32467_p3) + $signed(lhs_52_fu_35132_p3));

assign p_Val2_365_fu_36080_p2 = ($signed(rhs_62_fu_32615_p3) + $signed(lhs_53_fu_35234_p3));

assign p_Val2_367_fu_38407_p2 = ($signed(rhs_63_fu_36277_p3) + $signed(lhs_54_reg_42896));

assign p_Val2_369_fu_38507_p2 = ($signed(rhs_64_fu_36402_p3) + $signed(lhs_55_reg_42902));

assign p_Val2_36_fu_19583_p2 = ($signed(zext_ln377_12_fu_19580_p1) + $signed(sext_ln823_12_fu_19577_p1));

assign p_Val2_371_fu_38607_p2 = ($signed(rhs_65_fu_36527_p3) + $signed(lhs_56_reg_42908));

assign p_Val2_373_fu_38707_p2 = ($signed(rhs_66_fu_36652_p3) + $signed(lhs_57_reg_42914));

assign p_Val2_375_fu_38807_p2 = ($signed(rhs_67_fu_36777_p3) + $signed(lhs_58_reg_42920));

assign p_Val2_377_fu_38907_p2 = ($signed(rhs_68_fu_36795_p3) + $signed(lhs_59_reg_42926));

assign p_Val2_379_fu_39007_p2 = ($signed(rhs_69_fu_36919_p3) + $signed(lhs_60_reg_42932));

assign p_Val2_381_fu_39107_p2 = ($signed(rhs_70_fu_37044_p3) + $signed(lhs_61_reg_42938));

assign p_Val2_383_fu_39207_p2 = ($signed(rhs_71_fu_37169_p3) + $signed(lhs_62_reg_42944));

assign p_Val2_385_fu_39308_p2 = ($signed(rhs_72_fu_37318_p3) + $signed(lhs_63_fu_38478_p3));

assign p_Val2_387_fu_39410_p2 = ($signed(rhs_73_fu_37467_p3) + $signed(lhs_64_fu_38578_p3));

assign p_Val2_389_fu_39512_p2 = ($signed(rhs_74_fu_37616_p3) + $signed(lhs_65_fu_38678_p3));

assign p_Val2_391_fu_39614_p2 = ($signed(rhs_75_fu_37765_p3) + $signed(lhs_66_fu_38778_p3));

assign p_Val2_393_fu_39716_p2 = ($signed(rhs_76_fu_37783_p3) + $signed(lhs_67_fu_38878_p3));

assign p_Val2_395_fu_39818_p2 = ($signed(rhs_77_fu_37931_p3) + $signed(lhs_68_fu_38978_p3));

assign p_Val2_397_fu_39920_p2 = ($signed(rhs_78_fu_38080_p3) + $signed(lhs_69_fu_39078_p3));

assign p_Val2_399_fu_40022_p2 = ($signed(rhs_79_fu_38229_p3) + $signed(lhs_70_fu_39178_p3));

assign p_Val2_39_fu_19732_p2 = ($signed(zext_ln377_13_fu_19729_p1) + $signed(sext_ln823_13_fu_19726_p1));

assign p_Val2_401_fu_40124_p2 = ($signed(rhs_80_fu_38378_p3) + $signed(lhs_71_fu_39278_p3));

assign p_Val2_40_fu_17597_p1 = p_read1_int_reg;

assign p_Val2_40_fu_17597_p4 = {{p_Val2_40_fu_17597_p1[31:16]}};

assign p_Val2_41_fu_17631_p2 = ($signed(zext_ln377_14_fu_17627_p1) + $signed(sext_ln823_2_fu_17607_p1));

assign p_Val2_43_fu_17749_p4 = {{r_V_12_fu_489_p2[41:24]}};

assign p_Val2_44_fu_17783_p2 = ($signed(zext_ln377_15_fu_17779_p1) + $signed(sext_ln823_14_fu_17759_p1));

assign p_Val2_47_fu_20023_p2 = ($signed(zext_ln377_16_fu_20020_p1) + $signed(sext_ln823_15_fu_20017_p1));

assign p_Val2_4_fu_16355_p4 = {{r_V_1_fu_470_p2[41:24]}};

assign p_Val2_50_fu_20172_p2 = ($signed(zext_ln377_17_fu_20169_p1) + $signed(sext_ln823_16_fu_20166_p1));

assign p_Val2_53_fu_20321_p2 = ($signed(zext_ln377_18_fu_20318_p1) + $signed(sext_ln823_17_fu_20315_p1));

assign p_Val2_56_fu_20450_p2 = ($signed(zext_ln377_19_fu_20447_p1) + $signed(sext_ln823_18_fu_20444_p1));

assign p_Val2_59_fu_20579_p2 = ($signed(zext_ln377_20_fu_20576_p1) + $signed(sext_ln823_19_fu_20573_p1));

assign p_Val2_5_fu_16389_p2 = ($signed(zext_ln377_1_fu_16385_p1) + $signed(sext_ln823_4_fu_16365_p1));

assign p_Val2_62_fu_20728_p2 = ($signed(zext_ln377_21_fu_20725_p1) + $signed(sext_ln823_20_fu_20722_p1));

assign p_Val2_65_fu_20857_p2 = ($signed(zext_ln377_22_fu_20854_p1) + $signed(sext_ln823_21_fu_20851_p1));

assign p_Val2_68_fu_20986_p2 = ($signed(zext_ln377_23_fu_20983_p1) + $signed(sext_ln823_22_fu_20980_p1));

assign p_Val2_70_fu_18207_p4 = {{r_V_21_fu_18193_p2[38:24]}};

assign p_Val2_71_fu_18241_p2 = ($signed(zext_ln377_24_fu_18237_p1) + $signed(sext_ln823_23_fu_18217_p1));

assign p_Val2_74_fu_21132_p2 = ($signed(zext_ln377_25_fu_21129_p1) + $signed(sext_ln823_24_fu_21126_p1));

assign p_Val2_77_fu_21261_p2 = ($signed(zext_ln377_26_fu_21258_p1) + $signed(sext_ln823_25_fu_21255_p1));

assign p_Val2_79_fu_21416_p4 = {{r_V_24_fu_508_p2[55:24]}};

assign p_Val2_7_fu_16449_p4 = {{r_V_2_fu_16435_p2[38:24]}};

assign p_Val2_80_fu_21446_p2 = (zext_ln377_27_fu_21442_p1 + p_Val2_79_fu_21416_p4);

assign p_Val2_82_fu_21476_p4 = {{r_V_25_fu_497_p2[43:24]}};

assign p_Val2_83_fu_21510_p2 = ($signed(zext_ln377_28_fu_21506_p1) + $signed(sext_ln823_26_fu_21486_p1));

assign p_Val2_85_fu_21540_p4 = {{r_V_26_fu_490_p2[42:24]}};

assign p_Val2_86_fu_21574_p2 = ($signed(zext_ln377_29_fu_21570_p1) + $signed(sext_ln823_27_fu_21550_p1));

assign p_Val2_88_fu_21604_p4 = {{r_V_27_fu_541_p2[43:24]}};

assign p_Val2_89_fu_21638_p2 = ($signed(zext_ln377_30_fu_21634_p1) + $signed(sext_ln823_28_fu_21614_p1));

assign p_Val2_8_fu_16489_p2 = ($signed(zext_ln377_2_fu_16485_p1) + $signed(sext_ln823_5_fu_16459_p1));

assign p_Val2_91_fu_21668_p4 = {{r_V_28_fu_521_p2[42:24]}};

assign p_Val2_92_fu_21702_p2 = ($signed(zext_ln377_31_fu_21698_p1) + $signed(sext_ln823_29_fu_21678_p1));

assign p_Val2_94_fu_21732_p4 = {{r_V_29_fu_538_p2[40:24]}};

assign p_Val2_95_fu_21766_p2 = ($signed(zext_ln377_32_fu_21762_p1) + $signed(sext_ln823_30_fu_21742_p1));

assign p_Val2_97_fu_21796_p4 = {{r_V_30_fu_488_p2[40:24]}};

assign p_Val2_98_fu_21830_p2 = ($signed(zext_ln377_33_fu_21826_p1) + $signed(sext_ln823_31_fu_21806_p1));

assign r_V_10_fu_548_p0 = sext_ln70_7_fu_17134_p1;

assign r_V_10_fu_548_p1 = 45'd2984;

assign r_V_11_fu_478_p0 = sext_ln70_7_fu_17134_p1;

assign r_V_11_fu_478_p1 = 45'd35184372086172;

assign r_V_12_fu_489_p1 = 42'd4398046510823;

assign r_V_13_fu_501_p0 = sext_ln70_8_fu_17141_p1;

assign r_V_13_fu_501_p1 = 43'd8796093021547;

assign r_V_14_fu_546_p0 = sext_ln70_7_fu_17134_p1;

assign r_V_14_fu_546_p1 = 45'd2054;

assign r_V_15_fu_482_p0 = sext_ln70_13_fu_17909_p1;

assign r_V_15_fu_482_p1 = 43'd530;

assign r_V_16_fu_492_p1 = 44'd1352;

assign r_V_17_fu_485_p1 = 42'd433;

assign r_V_18_fu_481_p0 = sext_ln70_13_fu_17909_p1;

assign r_V_18_fu_481_p1 = 43'd8796093021244;

assign r_V_19_fu_473_p0 = sext_ln70_13_fu_17909_p1;

assign r_V_19_fu_473_p1 = 43'd999;

assign r_V_1_fu_470_p1 = 42'd266;

assign r_V_20_fu_515_p1 = 38'd274877906921;

assign r_V_21_fu_18193_p2 = ($signed(sext_ln1273_1_fu_18177_p1) - $signed(sext_ln1273_2_fu_18189_p1));

assign r_V_22_fu_535_p1 = 45'd35184372086441;

assign r_V_23_fu_518_p0 = sext_ln70_13_fu_17909_p1;

assign r_V_23_fu_518_p1 = 43'd8796093021444;

assign r_V_24_fu_508_p0 = sext_ln70_18_fu_21403_p1;

assign r_V_24_fu_508_p1 = 56'd10490509;

assign r_V_25_fu_497_p0 = sext_ln70_17_fu_21398_p1;

assign r_V_25_fu_497_p1 = 44'd17592186042933;

assign r_V_26_fu_490_p0 = sext_ln70_16_fu_21393_p1;

assign r_V_26_fu_490_p1 = 43'd566;

assign r_V_27_fu_541_p0 = sext_ln70_17_fu_21398_p1;

assign r_V_27_fu_541_p1 = 44'd17592186043385;

assign r_V_28_fu_521_p0 = sext_ln70_16_fu_21393_p1;

assign r_V_28_fu_521_p1 = 43'd819;

assign r_V_29_fu_538_p0 = sext_ln70_15_fu_21388_p1;

assign r_V_29_fu_538_p1 = 41'd2199023255329;

assign r_V_2_fu_16435_p2 = ($signed(sext_ln70_3_fu_16269_p1) - $signed(sext_ln1273_fu_16419_p1));

assign r_V_30_fu_488_p0 = sext_ln70_15_fu_21388_p1;

assign r_V_30_fu_488_p1 = 41'd2199023255394;

assign r_V_31_fu_496_p1 = 46'd70368744170099;

assign r_V_32_fu_499_p0 = sext_ln70_18_fu_21403_p1;

assign r_V_32_fu_499_p1 = 56'd72057594028989239;

assign r_V_33_fu_527_p1 = 51'd2251799813319069;

assign r_V_34_fu_509_p0 = sext_ln70_24_fu_21996_p1;

assign r_V_34_fu_509_p1 = 44'd17592186043320;

assign r_V_35_fu_476_p1 = 42'd291;

assign r_V_36_fu_22142_p2 = ($signed(sext_ln1273_3_fu_22138_p1) - $signed(sext_ln70_22_fu_21989_p1));

assign r_V_37_fu_494_p0 = sext_ln70_21_fu_21984_p1;

assign r_V_37_fu_494_p1 = 43'd639;

assign r_V_38_fu_498_p0 = sext_ln70_24_fu_21996_p1;

assign r_V_38_fu_498_p1 = 44'd17592186042810;

assign r_V_39_fu_505_p0 = sext_ln70_21_fu_21984_p1;

assign r_V_39_fu_505_p1 = 43'd8796093021539;

assign r_V_3_fu_510_p0 = sext_ln70_2_fu_16263_p1;

assign r_V_3_fu_510_p1 = 45'd35184372086226;

assign r_V_40_fu_512_p1 = 45'd3204;

assign r_V_41_fu_472_p1 = 53'd1562550;

assign r_V_42_fu_26887_p2 = ($signed(sext_ln70_30_fu_26873_p1) - $signed(sext_ln1273_4_fu_26883_p1));

assign r_V_43_fu_531_p0 = sext_ln70_29_fu_26867_p1;

assign r_V_43_fu_531_p1 = 43'd8796093021305;

assign r_V_44_fu_520_p1 = 42'd4398046510717;

assign r_V_45_fu_506_p1 = 45'd2399;

assign r_V_46_fu_530_p1 = 44'd17592186043315;

assign r_V_47_fu_471_p0 = sext_ln70_29_fu_26867_p1;

assign r_V_47_fu_471_p1 = 43'd657;

assign r_V_48_fu_27412_p2 = ($signed(sub_ln1273_fu_27395_p2) - $signed(sext_ln1273_6_fu_27408_p1));

assign r_V_49_fu_480_p0 = sext_ln70_29_fu_26867_p1;

assign r_V_49_fu_480_p1 = 43'd8796093021646;

assign r_V_4_fu_526_p0 = sext_ln70_1_fu_16257_p1;

assign r_V_4_fu_526_p1 = 43'd8796093021339;

assign r_V_50_fu_27673_p2 = ($signed(sext_ln1273_5_fu_27391_p1) - $signed(sext_ln1273_7_fu_27669_p1));

assign r_V_51_fu_491_p1 = 43'd615;

assign r_V_52_fu_523_p1 = 42'd4398046510611;

assign r_V_53_fu_534_p0 = sext_ln70_32_fu_27865_p1;

assign r_V_53_fu_534_p1 = 44'd1741;

assign r_V_54_fu_493_p0 = sext_ln70_31_fu_27859_p1;

assign r_V_54_fu_493_p1 = 45'd35184372085507;

assign r_V_55_fu_540_p0 = sext_ln70_31_fu_27859_p1;

assign r_V_55_fu_540_p1 = 45'd3186;

assign r_V_56_fu_549_p0 = sext_ln70_32_fu_27865_p1;

assign r_V_56_fu_549_p1 = 44'd17592186042977;

assign r_V_57_fu_504_p0 = sext_ln70_31_fu_27859_p1;

assign r_V_57_fu_504_p1 = 45'd35184372086664;

assign r_V_58_fu_28195_p2 = ($signed(sext_ln1273_8_fu_28180_p1) - $signed(sext_ln1273_9_fu_28191_p1));

assign r_V_59_fu_532_p0 = sext_ln70_32_fu_27865_p1;

assign r_V_59_fu_532_p1 = 44'd17592186043197;

assign r_V_5_fu_500_p0 = sext_ln70_1_fu_16257_p1;

assign r_V_5_fu_500_p1 = 43'd8796093021348;

assign r_V_60_fu_474_p0 = sext_ln70_37_fu_32634_p1;

assign r_V_60_fu_474_p1 = 42'd4398046510813;

assign r_V_61_fu_543_p0 = sext_ln70_36_fu_32629_p1;

assign r_V_61_fu_543_p1 = 43'd970;

assign r_V_62_fu_477_p0 = sext_ln70_35_fu_32623_p1;

assign r_V_62_fu_477_p1 = 44'd1347;

assign r_V_63_fu_545_p0 = sext_ln70_37_fu_32634_p1;

assign r_V_63_fu_545_p1 = 42'd4398046510679;

assign r_V_64_fu_533_p0 = sext_ln70_35_fu_32623_p1;

assign r_V_64_fu_533_p1 = 44'd1766;

assign r_V_65_fu_32971_p2 = ($signed(39'd0) - $signed(sext_ln1273_10_fu_32967_p1));

assign r_V_66_fu_511_p0 = sext_ln70_36_fu_32629_p1;

assign r_V_66_fu_511_p1 = 43'd8796093021501;

assign r_V_67_fu_522_p0 = sext_ln70_35_fu_32623_p1;

assign r_V_67_fu_522_p1 = 44'd17592186043389;

assign r_V_68_fu_544_p0 = sext_ln70_37_fu_32634_p1;

assign r_V_68_fu_544_p1 = 42'd4398046510785;

assign r_V_69_fu_529_p1 = 44'd17592186043131;

assign r_V_6_fu_16819_p2 = ($signed(39'd0) - $signed(sext_ln1273_fu_16419_p1));

assign r_V_70_fu_516_p0 = sext_ln70_43_fu_33369_p1;

assign r_V_70_fu_516_p1 = 43'd547;

assign r_V_71_fu_517_p1 = 42'd4398046510692;

assign r_V_72_fu_525_p0 = sext_ln70_43_fu_33369_p1;

assign r_V_72_fu_525_p1 = 43'd8796093021555;

assign r_V_73_fu_33568_p2 = ($signed(sext_ln1273_11_fu_33553_p1) - $signed(sext_ln1273_12_fu_33564_p1));

assign r_V_74_fu_495_p1 = 41'd2199023255382;

assign r_V_75_fu_539_p1 = 40'd125;

assign r_V_76_fu_484_p1 = 46'd5882;

assign r_V_77_fu_486_p1 = 54'd3281710;

assign r_V_7_fu_537_p1 = 57'd144115188051572030;

assign r_V_8_fu_514_p0 = sext_ln70_2_fu_16263_p1;

assign r_V_8_fu_514_p1 = 45'd3212;

assign r_V_9_fu_503_p0 = sext_ln70_8_fu_17141_p1;

assign r_V_9_fu_503_p1 = 43'd529;

assign r_V_fu_519_p1 = 47'd140737488340165;

assign ret_V_10_fu_23530_p2 = ($signed(sext_ln813_12_fu_23526_p1) + $signed(sext_ln813_11_fu_23522_p1));

assign ret_V_11_fu_23632_p2 = ($signed(sext_ln813_14_fu_23628_p1) + $signed(sext_ln813_13_fu_23624_p1));

assign ret_V_12_fu_23734_p2 = ($signed(sext_ln813_16_fu_23730_p1) + $signed(sext_ln813_15_fu_23726_p1));

assign ret_V_13_fu_23836_p2 = ($signed(sext_ln813_18_fu_23832_p1) + $signed(sext_ln813_17_fu_23828_p1));

assign ret_V_14_fu_23938_p2 = ($signed(sext_ln813_20_fu_23934_p1) + $signed(sext_ln813_19_fu_23930_p1));

assign ret_V_15_fu_24040_p2 = ($signed(sext_ln813_22_fu_24036_p1) + $signed(sext_ln813_21_fu_24032_p1));

assign ret_V_16_fu_24142_p2 = ($signed(sext_ln813_24_fu_24138_p1) + $signed(sext_ln813_23_fu_24134_p1));

assign ret_V_17_fu_24244_p2 = ($signed(sext_ln813_26_fu_24240_p1) + $signed(sext_ln813_25_fu_24236_p1));

assign ret_V_18_fu_28430_p2 = ($signed(sext_ln813_28_fu_28426_p1) + $signed(sext_ln813_27_fu_28423_p1));

assign ret_V_19_fu_28530_p2 = ($signed(sext_ln813_30_fu_28526_p1) + $signed(sext_ln813_29_fu_28523_p1));

assign ret_V_1_fu_22640_p2 = ($signed(sext_ln813_1_fu_22636_p1) + $signed(33'd8589738296));

assign ret_V_20_fu_24346_p2 = ($signed(sext_ln813_32_fu_24342_p1) + $signed(sext_ln813_31_fu_24338_p1));

assign ret_V_21_fu_28688_p2 = ($signed(sext_ln813_34_fu_28684_p1) + $signed(sext_ln813_33_fu_28681_p1));

assign ret_V_22_fu_28788_p2 = ($signed(sext_ln813_36_fu_28784_p1) + $signed(sext_ln813_35_fu_28781_p1));

assign ret_V_23_fu_28888_p2 = ($signed(sext_ln813_38_fu_28884_p1) + $signed(sext_ln813_37_fu_28881_p1));

assign ret_V_24_fu_24382_p2 = ($signed(sext_ln813_40_fu_24378_p1) + $signed(sext_ln813_39_fu_24374_p1));

assign ret_V_25_fu_29046_p2 = ($signed(sext_ln813_42_fu_29042_p1) + $signed(sext_ln813_41_fu_29039_p1));

assign ret_V_26_fu_29146_p2 = ($signed(sext_ln813_44_fu_29142_p1) + $signed(sext_ln813_43_fu_29139_p1));

assign ret_V_27_fu_29247_p2 = ($signed(sext_ln813_46_fu_29243_p1) + $signed(sext_ln813_45_fu_29239_p1));

assign ret_V_28_fu_29349_p2 = ($signed(sext_ln813_48_fu_29345_p1) + $signed(sext_ln813_47_fu_29341_p1));

assign ret_V_29_fu_29451_p2 = ($signed(sext_ln813_50_fu_29447_p1) + $signed(sext_ln813_49_fu_29443_p1));

assign ret_V_2_fu_22738_p2 = ($signed(sext_ln813_2_fu_22734_p1) + $signed(33'd8588322428));

assign ret_V_30_fu_29553_p2 = ($signed(sext_ln813_52_fu_29549_p1) + $signed(sext_ln813_51_fu_29545_p1));

assign ret_V_31_fu_29655_p2 = ($signed(sext_ln813_54_fu_29651_p1) + $signed(sext_ln813_53_fu_29647_p1));

assign ret_V_32_fu_29757_p2 = ($signed(sext_ln813_56_fu_29753_p1) + $signed(sext_ln813_55_fu_29749_p1));

assign ret_V_33_fu_29859_p2 = ($signed(sext_ln813_58_fu_29855_p1) + $signed(sext_ln813_57_fu_29851_p1));

assign ret_V_34_fu_29961_p2 = ($signed(sext_ln813_60_fu_29957_p1) + $signed(sext_ln813_59_fu_29953_p1));

assign ret_V_35_fu_30063_p2 = ($signed(sext_ln813_62_fu_30059_p1) + $signed(sext_ln813_61_fu_30055_p1));

assign ret_V_36_fu_30165_p2 = ($signed(sext_ln813_64_fu_30161_p1) + $signed(sext_ln813_63_fu_30157_p1));

assign ret_V_37_fu_30201_p2 = ($signed(sext_ln813_66_fu_30197_p1) + $signed(sext_ln813_65_fu_30193_p1));

assign ret_V_38_fu_30237_p2 = ($signed(sext_ln813_68_fu_30233_p1) + $signed(sext_ln813_67_fu_30229_p1));

assign ret_V_39_fu_30339_p2 = ($signed(sext_ln813_70_fu_30335_p1) + $signed(sext_ln813_69_fu_30331_p1));

assign ret_V_3_fu_22836_p2 = ($signed(sext_ln813_3_fu_22832_p1) + $signed(33'd8588872678));

assign ret_V_40_fu_30375_p2 = ($signed(sext_ln813_72_fu_30371_p1) + $signed(sext_ln813_71_fu_30367_p1));

assign ret_V_41_fu_30411_p2 = ($signed(sext_ln813_74_fu_30407_p1) + $signed(sext_ln813_73_fu_30403_p1));

assign ret_V_42_fu_30447_p2 = ($signed(sext_ln813_76_fu_30443_p1) + $signed(sext_ln813_75_fu_30439_p1));

assign ret_V_43_fu_30549_p2 = ($signed(sext_ln813_78_fu_30545_p1) + $signed(sext_ln813_77_fu_30541_p1));

assign ret_V_44_fu_30585_p2 = ($signed(sext_ln813_80_fu_30581_p1) + $signed(sext_ln813_79_fu_30577_p1));

assign ret_V_45_fu_34336_p2 = ($signed(sext_ln813_82_fu_34332_p1) + $signed(sext_ln813_81_fu_34328_p1));

assign ret_V_46_fu_34438_p2 = ($signed(sext_ln813_84_fu_34434_p1) + $signed(sext_ln813_83_fu_34430_p1));

assign ret_V_47_fu_34539_p2 = ($signed(sext_ln813_86_fu_34535_p1) + $signed(sext_ln813_85_fu_34532_p1));

assign ret_V_48_fu_34640_p2 = ($signed(sext_ln813_88_fu_34636_p1) + $signed(sext_ln813_87_fu_34632_p1));

assign ret_V_49_fu_34742_p2 = ($signed(sext_ln813_90_fu_34738_p1) + $signed(sext_ln813_89_fu_34734_p1));

assign ret_V_4_fu_22934_p2 = ($signed(sext_ln813_4_fu_22930_p1) + $signed(33'd8589930257));

assign ret_V_50_fu_34844_p2 = ($signed(sext_ln813_92_fu_34840_p1) + $signed(sext_ln813_91_fu_34836_p1));

assign ret_V_51_fu_34945_p2 = ($signed(sext_ln813_94_fu_34941_p1) + $signed(sext_ln813_93_fu_34938_p1));

assign ret_V_52_fu_35046_p2 = ($signed(sext_ln813_96_fu_35042_p1) + $signed(sext_ln813_95_fu_35038_p1));

assign ret_V_53_fu_35148_p2 = ($signed(sext_ln813_98_fu_35144_p1) + $signed(sext_ln813_97_fu_35140_p1));

assign ret_V_54_fu_35250_p2 = ($signed(sext_ln813_100_fu_35246_p1) + $signed(sext_ln813_99_fu_35242_p1));

assign ret_V_55_fu_35352_p2 = ($signed(sext_ln813_102_fu_35348_p1) + $signed(sext_ln813_101_fu_35344_p1));

assign ret_V_56_fu_35454_p2 = ($signed(sext_ln813_104_fu_35450_p1) + $signed(sext_ln813_103_fu_35446_p1));

assign ret_V_57_fu_35556_p2 = ($signed(sext_ln813_106_fu_35552_p1) + $signed(sext_ln813_105_fu_35548_p1));

assign ret_V_58_fu_35658_p2 = ($signed(sext_ln813_108_fu_35654_p1) + $signed(sext_ln813_107_fu_35650_p1));

assign ret_V_59_fu_35760_p2 = ($signed(sext_ln813_110_fu_35756_p1) + $signed(sext_ln813_109_fu_35752_p1));

assign ret_V_5_fu_23032_p2 = ($signed(sext_ln813_5_fu_23028_p1) + $signed(33'd8589928913));

assign ret_V_60_fu_35862_p2 = ($signed(sext_ln813_112_fu_35858_p1) + $signed(sext_ln813_111_fu_35854_p1));

assign ret_V_61_fu_35964_p2 = ($signed(sext_ln813_114_fu_35960_p1) + $signed(sext_ln813_113_fu_35956_p1));

assign ret_V_62_fu_36066_p2 = ($signed(sext_ln813_116_fu_36062_p1) + $signed(sext_ln813_115_fu_36058_p1));

assign ret_V_63_fu_38393_p2 = ($signed(sext_ln813_118_fu_38389_p1) + $signed(sext_ln813_117_fu_38386_p1));

assign ret_V_64_fu_38493_p2 = ($signed(sext_ln813_120_fu_38489_p1) + $signed(sext_ln813_119_fu_38486_p1));

assign ret_V_65_fu_38593_p2 = ($signed(sext_ln813_122_fu_38589_p1) + $signed(sext_ln813_121_fu_38586_p1));

assign ret_V_66_fu_38693_p2 = ($signed(sext_ln813_124_fu_38689_p1) + $signed(sext_ln813_123_fu_38686_p1));

assign ret_V_67_fu_38793_p2 = ($signed(sext_ln813_126_fu_38789_p1) + $signed(sext_ln813_125_fu_38786_p1));

assign ret_V_68_fu_38893_p2 = ($signed(sext_ln813_128_fu_38889_p1) + $signed(sext_ln813_127_fu_38886_p1));

assign ret_V_69_fu_38993_p2 = ($signed(sext_ln813_130_fu_38989_p1) + $signed(sext_ln813_129_fu_38986_p1));

assign ret_V_6_fu_23130_p2 = ($signed(sext_ln813_6_fu_23126_p1) + $signed(33'd8589908017));

assign ret_V_70_fu_39093_p2 = ($signed(sext_ln813_132_fu_39089_p1) + $signed(sext_ln813_131_fu_39086_p1));

assign ret_V_71_fu_39193_p2 = ($signed(sext_ln813_134_fu_39189_p1) + $signed(sext_ln813_133_fu_39186_p1));

assign ret_V_72_fu_39294_p2 = ($signed(sext_ln813_136_fu_39290_p1) + $signed(sext_ln813_135_fu_39286_p1));

assign ret_V_73_fu_39396_p2 = ($signed(sext_ln813_138_fu_39392_p1) + $signed(sext_ln813_137_fu_39388_p1));

assign ret_V_74_fu_39498_p2 = ($signed(sext_ln813_140_fu_39494_p1) + $signed(sext_ln813_139_fu_39490_p1));

assign ret_V_75_fu_39600_p2 = ($signed(sext_ln813_142_fu_39596_p1) + $signed(sext_ln813_141_fu_39592_p1));

assign ret_V_76_fu_39702_p2 = ($signed(sext_ln813_144_fu_39698_p1) + $signed(sext_ln813_143_fu_39694_p1));

assign ret_V_77_fu_39804_p2 = ($signed(sext_ln813_146_fu_39800_p1) + $signed(sext_ln813_145_fu_39796_p1));

assign ret_V_78_fu_39906_p2 = ($signed(sext_ln813_148_fu_39902_p1) + $signed(sext_ln813_147_fu_39898_p1));

assign ret_V_79_fu_40008_p2 = ($signed(sext_ln813_150_fu_40004_p1) + $signed(sext_ln813_149_fu_40000_p1));

assign ret_V_7_fu_23228_p2 = ($signed(sext_ln813_7_fu_23224_p1) + $signed(33'd5062185));

assign ret_V_80_fu_40110_p2 = ($signed(sext_ln813_152_fu_40106_p1) + $signed(sext_ln813_151_fu_40102_p1));

assign ret_V_8_fu_23326_p2 = ($signed(sext_ln813_8_fu_23322_p1) + $signed(33'd6923874));

assign ret_V_9_fu_23428_p2 = ($signed(sext_ln813_10_fu_23424_p1) + $signed(sext_ln813_9_fu_23420_p1));

assign ret_V_fu_22542_p2 = ($signed(sext_ln813_fu_22538_p1) + $signed(33'd140968));

assign rhs_10_fu_19553_p3 = ((or_ln346_10_reg_40609[0:0] == 1'b1) ? select_ln346_20_fu_19546_p3 : sext_ln856_fu_19543_p1);

assign rhs_11_fu_19570_p3 = ((or_ln346_11_reg_40624[0:0] == 1'b1) ? select_ln346_22_fu_19563_p3 : sext_ln856_1_fu_19560_p1);

assign rhs_12_fu_19718_p3 = ((or_ln346_12_fu_19712_p2[0:0] == 1'b1) ? select_ln346_24_fu_19704_p3 : sext_ln856_12_fu_19589_p1);

assign rhs_13_fu_19867_p3 = ((or_ln346_13_fu_19861_p2[0:0] == 1'b1) ? select_ln346_26_fu_19853_p3 : sext_ln856_13_fu_19738_p1);

assign rhs_14_fu_19885_p3 = ((or_ln346_14_reg_40697[0:0] == 1'b1) ? select_ln346_28_fu_19878_p3 : sext_ln856_2_fu_19875_p1);

assign rhs_15_fu_20009_p3 = ((or_ln346_15_fu_20003_p2[0:0] == 1'b1) ? select_ln346_30_fu_19995_p3 : sext_ln856_14_fu_19892_p1);

assign rhs_16_fu_20158_p3 = ((or_ln346_16_fu_20152_p2[0:0] == 1'b1) ? select_ln346_32_fu_20144_p3 : sext_ln856_15_fu_20029_p1);

assign rhs_17_fu_20307_p3 = ((or_ln346_17_fu_20301_p2[0:0] == 1'b1) ? select_ln346_34_fu_20293_p3 : sext_ln856_16_fu_20178_p1);

assign rhs_18_fu_24420_p3 = ((or_ln346_18_reg_41053[0:0] == 1'b1) ? select_ln346_36_fu_24413_p3 : sext_ln856_17_fu_24410_p1);

assign rhs_19_fu_24437_p3 = ((or_ln346_19_reg_41068[0:0] == 1'b1) ? select_ln346_38_fu_24430_p3 : sext_ln856_18_fu_24427_p1);

assign rhs_1_fu_18731_p3 = ((or_ln346_1_fu_18725_p2[0:0] == 1'b1) ? select_ln346_2_fu_18717_p3 : sext_ln856_4_fu_18614_p1);

assign rhs_20_fu_20714_p3 = ((or_ln346_20_fu_20708_p2[0:0] == 1'b1) ? select_ln346_40_fu_20700_p3 : sext_ln856_19_fu_20585_p1);

assign rhs_21_fu_24454_p3 = ((or_ln346_21_reg_41083[0:0] == 1'b1) ? select_ln346_42_fu_24447_p3 : sext_ln856_20_fu_24444_p1);

assign rhs_22_fu_24471_p3 = ((or_ln346_22_reg_41098[0:0] == 1'b1) ? select_ln346_44_fu_24464_p3 : sext_ln856_21_fu_24461_p1);

assign rhs_23_fu_24488_p3 = ((or_ln346_23_reg_41113[0:0] == 1'b1) ? select_ln346_46_fu_24481_p3 : sext_ln856_22_fu_24478_p1);

assign rhs_24_fu_21119_p3 = ((or_ln346_24_reg_40975[0:0] == 1'b1) ? select_ln346_48_fu_21112_p3 : sext_ln856_23_fu_21109_p1);

assign rhs_25_fu_24505_p3 = ((or_ln346_25_reg_41128[0:0] == 1'b1) ? select_ln346_50_fu_24498_p3 : sext_ln856_24_fu_24495_p1);

assign rhs_26_fu_24522_p3 = ((or_ln346_26_reg_41143[0:0] == 1'b1) ? select_ln346_52_fu_24515_p3 : sext_ln856_25_fu_24512_p1);

assign rhs_27_fu_24643_p3 = ((or_ln346_27_fu_24637_p2[0:0] == 1'b1) ? select_ln346_54_fu_24629_p3 : p_Val2_80_reg_41160);

assign rhs_28_fu_24767_p3 = ((or_ln346_28_fu_24761_p2[0:0] == 1'b1) ? select_ln346_56_fu_24753_p3 : sext_ln856_26_fu_24650_p1);

assign rhs_29_fu_24892_p3 = ((or_ln346_29_fu_24886_p2[0:0] == 1'b1) ? select_ln346_58_fu_24878_p3 : sext_ln856_27_fu_24775_p1);

assign rhs_2_fu_18749_p3 = ((or_ln346_2_reg_40395[0:0] == 1'b1) ? select_ln346_4_fu_18742_p3 : sext_ln856_5_fu_18739_p1);

assign rhs_30_fu_25017_p3 = ((or_ln346_30_fu_25011_p2[0:0] == 1'b1) ? select_ln346_60_fu_25003_p3 : sext_ln856_28_fu_24900_p1);

assign rhs_31_fu_25142_p3 = ((or_ln346_31_fu_25136_p2[0:0] == 1'b1) ? select_ln346_62_fu_25128_p3 : sext_ln856_29_fu_25025_p1);

assign rhs_32_fu_25267_p3 = ((or_ln346_32_fu_25261_p2[0:0] == 1'b1) ? select_ln346_64_fu_25253_p3 : sext_ln856_30_fu_25150_p1);

assign rhs_33_fu_25392_p3 = ((or_ln346_33_fu_25386_p2[0:0] == 1'b1) ? select_ln346_66_fu_25378_p3 : sext_ln856_31_fu_25275_p1);

assign rhs_34_fu_25517_p3 = ((or_ln346_34_fu_25511_p2[0:0] == 1'b1) ? select_ln346_68_fu_25503_p3 : sext_ln856_32_fu_25400_p1);

assign rhs_35_fu_25639_p3 = ((or_ln346_35_fu_25633_p2[0:0] == 1'b1) ? select_ln346_70_fu_25625_p3 : p_Val2_104_reg_41408);

assign rhs_36_fu_25787_p3 = ((or_ln346_36_fu_25781_p2[0:0] == 1'b1) ? select_ln346_72_fu_25773_p3 : sext_ln856_33_fu_25658_p1);

assign rhs_37_fu_25936_p3 = ((or_ln346_37_fu_25930_p2[0:0] == 1'b1) ? select_ln346_74_fu_25922_p3 : sext_ln856_34_fu_25807_p1);

assign rhs_38_fu_26085_p3 = ((or_ln346_38_fu_26079_p2[0:0] == 1'b1) ? select_ln346_76_fu_26071_p3 : sext_ln856_35_fu_25956_p1);

assign rhs_39_fu_26103_p3 = ((or_ln346_39_reg_41524[0:0] == 1'b1) ? select_ln346_78_fu_26096_p3 : sext_ln856_36_fu_26093_p1);

assign rhs_3_fu_18873_p3 = ((or_ln346_3_fu_18867_p2[0:0] == 1'b1) ? select_ln346_6_fu_18859_p3 : sext_ln856_6_fu_18756_p1);

assign rhs_40_fu_26251_p3 = ((or_ln346_40_fu_26245_p2[0:0] == 1'b1) ? select_ln346_80_fu_26237_p3 : sext_ln856_37_fu_26122_p1);

assign rhs_41_fu_26400_p3 = ((or_ln346_41_fu_26394_p2[0:0] == 1'b1) ? select_ln346_82_fu_26386_p3 : sext_ln856_38_fu_26271_p1);

assign rhs_42_fu_26549_p3 = ((or_ln346_42_fu_26543_p2[0:0] == 1'b1) ? select_ln346_84_fu_26535_p3 : sext_ln856_39_fu_26420_p1);

assign rhs_43_fu_26698_p3 = ((or_ln346_43_fu_26692_p2[0:0] == 1'b1) ? select_ln346_86_fu_26684_p3 : sext_ln856_40_fu_26569_p1);

assign rhs_44_fu_26847_p3 = ((or_ln346_44_fu_26841_p2[0:0] == 1'b1) ? select_ln346_88_fu_26833_p3 : sext_ln856_41_fu_26718_p1);

assign rhs_45_fu_30623_p3 = ((or_ln346_45_reg_41766[0:0] == 1'b1) ? select_ln346_90_fu_30616_p3 : sext_ln856_42_fu_30613_p1);

assign rhs_46_fu_30747_p3 = ((or_ln346_46_fu_30741_p2[0:0] == 1'b1) ? select_ln346_92_fu_30733_p3 : sext_ln856_43_fu_30630_p1);

assign rhs_47_fu_30872_p3 = ((or_ln346_47_fu_30866_p2[0:0] == 1'b1) ? select_ln346_94_fu_30858_p3 : sext_ln856_44_fu_30755_p1);

assign rhs_48_fu_30997_p3 = ((or_ln346_48_fu_30991_p2[0:0] == 1'b1) ? select_ln346_96_fu_30983_p3 : sext_ln856_45_fu_30880_p1);

assign rhs_49_fu_31122_p3 = ((or_ln346_49_fu_31116_p2[0:0] == 1'b1) ? select_ln346_98_fu_31108_p3 : sext_ln856_46_fu_31005_p1);

assign rhs_4_fu_18998_p3 = ((or_ln346_4_fu_18992_p2[0:0] == 1'b1) ? select_ln346_8_fu_18984_p3 : sext_ln856_7_fu_18881_p1);

assign rhs_50_fu_31247_p3 = ((or_ln346_50_fu_31241_p2[0:0] == 1'b1) ? select_ln346_100_fu_31233_p3 : sext_ln856_47_fu_31130_p1);

assign rhs_51_fu_31265_p3 = ((or_ln346_51_reg_41936[0:0] == 1'b1) ? select_ln346_102_fu_31258_p3 : sext_ln856_48_fu_31255_p1);

assign rhs_52_fu_31389_p3 = ((or_ln346_52_fu_31383_p2[0:0] == 1'b1) ? select_ln346_104_fu_31375_p3 : sext_ln856_49_fu_31272_p1);

assign rhs_53_fu_31407_p3 = ((or_ln346_53_reg_41982[0:0] == 1'b1) ? select_ln346_106_fu_31400_p3 : sext_ln856_50_fu_31397_p1);

assign rhs_54_fu_31555_p3 = ((or_ln346_54_fu_31549_p2[0:0] == 1'b1) ? select_ln346_108_fu_31541_p3 : sext_ln856_51_fu_31426_p1);

assign rhs_55_fu_31704_p3 = ((or_ln346_55_fu_31698_p2[0:0] == 1'b1) ? select_ln346_110_fu_31690_p3 : sext_ln856_52_fu_31575_p1);

assign rhs_56_fu_31853_p3 = ((or_ln346_56_fu_31847_p2[0:0] == 1'b1) ? select_ln346_112_fu_31839_p3 : sext_ln856_53_fu_31724_p1);

assign rhs_57_fu_32002_p3 = ((or_ln346_57_fu_31996_p2[0:0] == 1'b1) ? select_ln346_114_fu_31988_p3 : sext_ln856_54_fu_31873_p1);

assign rhs_58_fu_32151_p3 = ((or_ln346_58_fu_32145_p2[0:0] == 1'b1) ? select_ln346_116_fu_32137_p3 : sext_ln856_55_fu_32022_p1);

assign rhs_59_fu_32300_p3 = ((or_ln346_59_fu_32294_p2[0:0] == 1'b1) ? select_ln346_118_fu_32286_p3 : sext_ln856_56_fu_32171_p1);

assign rhs_5_fu_19123_p3 = ((or_ln346_5_fu_19117_p2[0:0] == 1'b1) ? select_ln346_10_fu_19109_p3 : sext_ln856_8_fu_19006_p1);

assign rhs_60_fu_32449_p3 = ((or_ln346_60_fu_32443_p2[0:0] == 1'b1) ? select_ln346_120_fu_32435_p3 : sext_ln856_57_fu_32320_p1);

assign rhs_61_fu_32467_p3 = ((or_ln346_61_reg_42200[0:0] == 1'b1) ? select_ln346_122_fu_32460_p3 : sext_ln856_58_fu_32457_p1);

assign rhs_62_fu_32615_p3 = ((or_ln346_62_fu_32609_p2[0:0] == 1'b1) ? select_ln346_124_fu_32601_p3 : sext_ln856_59_fu_32486_p1);

assign rhs_63_fu_36277_p3 = ((or_ln346_63_fu_36271_p2[0:0] == 1'b1) ? select_ln346_126_fu_36263_p3 : sext_ln856_60_fu_36160_p1);

assign rhs_64_fu_36402_p3 = ((or_ln346_64_fu_36396_p2[0:0] == 1'b1) ? select_ln346_128_fu_36388_p3 : sext_ln856_61_fu_36285_p1);

assign rhs_65_fu_36527_p3 = ((or_ln346_65_fu_36521_p2[0:0] == 1'b1) ? select_ln346_130_fu_36513_p3 : sext_ln856_62_fu_36410_p1);

assign rhs_66_fu_36652_p3 = ((or_ln346_66_fu_36646_p2[0:0] == 1'b1) ? select_ln346_132_fu_36638_p3 : sext_ln856_63_fu_36535_p1);

assign rhs_67_fu_36777_p3 = ((or_ln346_67_fu_36771_p2[0:0] == 1'b1) ? select_ln346_134_fu_36763_p3 : sext_ln856_64_fu_36660_p1);

assign rhs_68_fu_36795_p3 = ((or_ln346_68_reg_42551[0:0] == 1'b1) ? select_ln346_136_fu_36788_p3 : sext_ln856_65_fu_36785_p1);

assign rhs_69_fu_36919_p3 = ((or_ln346_69_fu_36913_p2[0:0] == 1'b1) ? select_ln346_138_fu_36905_p3 : sext_ln856_66_fu_36802_p1);

assign rhs_6_fu_19141_p3 = ((or_ln346_6_reg_40503[0:0] == 1'b1) ? select_ln346_12_fu_19134_p3 : sext_ln856_9_fu_19131_p1);

assign rhs_70_fu_37044_p3 = ((or_ln346_70_fu_37038_p2[0:0] == 1'b1) ? select_ln346_140_fu_37030_p3 : sext_ln856_67_fu_36927_p1);

assign rhs_71_fu_37169_p3 = ((or_ln346_71_fu_37163_p2[0:0] == 1'b1) ? select_ln346_142_fu_37155_p3 : sext_ln856_68_fu_37052_p1);

assign rhs_72_fu_37318_p3 = ((or_ln346_72_fu_37312_p2[0:0] == 1'b1) ? select_ln346_144_fu_37304_p3 : sext_ln856_69_fu_37189_p1);

assign rhs_73_fu_37467_p3 = ((or_ln346_73_fu_37461_p2[0:0] == 1'b1) ? select_ln346_146_fu_37453_p3 : sext_ln856_70_fu_37338_p1);

assign rhs_74_fu_37616_p3 = ((or_ln346_74_fu_37610_p2[0:0] == 1'b1) ? select_ln346_148_fu_37602_p3 : sext_ln856_71_fu_37487_p1);

assign rhs_75_fu_37765_p3 = ((or_ln346_75_fu_37759_p2[0:0] == 1'b1) ? select_ln346_150_fu_37751_p3 : sext_ln856_72_fu_37636_p1);

assign rhs_76_fu_37783_p3 = ((or_ln346_76_reg_42775[0:0] == 1'b1) ? select_ln346_152_fu_37776_p3 : sext_ln856_73_fu_37773_p1);

assign rhs_77_fu_37931_p3 = ((or_ln346_77_fu_37925_p2[0:0] == 1'b1) ? select_ln346_154_fu_37917_p3 : sext_ln856_74_fu_37802_p1);

assign rhs_78_fu_38080_p3 = ((or_ln346_78_fu_38074_p2[0:0] == 1'b1) ? select_ln346_156_fu_38066_p3 : sext_ln856_75_fu_37951_p1);

assign rhs_79_fu_38229_p3 = ((or_ln346_79_fu_38223_p2[0:0] == 1'b1) ? select_ln346_158_fu_38215_p3 : sext_ln856_76_fu_38100_p1);

assign rhs_7_fu_19262_p3 = ((or_ln346_7_fu_19256_p2[0:0] == 1'b1) ? select_ln346_14_fu_19248_p3 : p_Val2_23_reg_40520);

assign rhs_80_fu_38378_p3 = ((or_ln346_80_fu_38372_p2[0:0] == 1'b1) ? select_ln346_160_fu_38364_p3 : sext_ln856_77_fu_38249_p1);

assign rhs_8_fu_19386_p3 = ((or_ln346_8_fu_19380_p2[0:0] == 1'b1) ? select_ln346_16_fu_19372_p3 : sext_ln856_10_fu_19269_p1);

assign rhs_9_fu_19535_p3 = ((or_ln346_9_fu_19529_p2[0:0] == 1'b1) ? select_ln346_18_fu_19521_p3 : sext_ln856_11_fu_19406_p1);

assign rhs_fu_18606_p3 = ((or_ln346_fu_18600_p2[0:0] == 1'b1) ? select_ln346_fu_18592_p3 : sext_ln856_3_fu_18489_p1);

assign select_ln302_100_fu_34914_p3 = ((xor_ln302_100_fu_34896_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_341_fu_34858_p2);

assign select_ln302_102_fu_35014_p3 = ((xor_ln302_102_fu_34996_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_343_fu_34959_p2);

assign select_ln302_104_fu_35116_p3 = ((xor_ln302_104_fu_35098_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_345_fu_35060_p2);

assign select_ln302_106_fu_35218_p3 = ((xor_ln302_106_fu_35200_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_347_fu_35162_p2);

assign select_ln302_108_fu_35320_p3 = ((xor_ln302_108_fu_35302_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_349_fu_35264_p2);

assign select_ln302_10_fu_23102_p3 = ((xor_ln302_10_fu_23084_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_251_fu_23046_p2);

assign select_ln302_110_fu_35422_p3 = ((xor_ln302_110_fu_35404_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_351_fu_35366_p2);

assign select_ln302_112_fu_35524_p3 = ((xor_ln302_112_fu_35506_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_353_fu_35468_p2);

assign select_ln302_114_fu_35626_p3 = ((xor_ln302_114_fu_35608_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_355_fu_35570_p2);

assign select_ln302_116_fu_35728_p3 = ((xor_ln302_116_fu_35710_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_357_fu_35672_p2);

assign select_ln302_118_fu_35830_p3 = ((xor_ln302_118_fu_35812_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_359_fu_35774_p2);

assign select_ln302_120_fu_35932_p3 = ((xor_ln302_120_fu_35914_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_361_fu_35876_p2);

assign select_ln302_122_fu_36034_p3 = ((xor_ln302_122_fu_36016_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_363_fu_35978_p2);

assign select_ln302_124_fu_36136_p3 = ((xor_ln302_124_fu_36118_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_365_fu_36080_p2);

assign select_ln302_126_fu_38462_p3 = ((xor_ln302_126_fu_38444_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_367_fu_38407_p2);

assign select_ln302_128_fu_38562_p3 = ((xor_ln302_128_fu_38544_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_369_fu_38507_p2);

assign select_ln302_12_fu_23200_p3 = ((xor_ln302_12_fu_23182_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_253_fu_23144_p2);

assign select_ln302_130_fu_38662_p3 = ((xor_ln302_130_fu_38644_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_371_fu_38607_p2);

assign select_ln302_132_fu_38762_p3 = ((xor_ln302_132_fu_38744_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_373_fu_38707_p2);

assign select_ln302_134_fu_38862_p3 = ((xor_ln302_134_fu_38844_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_375_fu_38807_p2);

assign select_ln302_136_fu_38962_p3 = ((xor_ln302_136_fu_38944_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_377_fu_38907_p2);

assign select_ln302_138_fu_39062_p3 = ((xor_ln302_138_fu_39044_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_379_fu_39007_p2);

assign select_ln302_140_fu_39162_p3 = ((xor_ln302_140_fu_39144_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_381_fu_39107_p2);

assign select_ln302_142_fu_39262_p3 = ((xor_ln302_142_fu_39244_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_383_fu_39207_p2);

assign select_ln302_144_fu_39364_p3 = ((xor_ln302_144_fu_39346_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_385_fu_39308_p2);

assign select_ln302_145_fu_39380_p3 = ((or_ln302_72_fu_39358_p2[0:0] == 1'b1) ? select_ln302_144_fu_39364_p3 : select_ln350_72_fu_39372_p3);

assign select_ln302_146_fu_39466_p3 = ((xor_ln302_146_fu_39448_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_387_fu_39410_p2);

assign select_ln302_147_fu_39482_p3 = ((or_ln302_73_fu_39460_p2[0:0] == 1'b1) ? select_ln302_146_fu_39466_p3 : select_ln350_73_fu_39474_p3);

assign select_ln302_148_fu_39568_p3 = ((xor_ln302_148_fu_39550_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_389_fu_39512_p2);

assign select_ln302_149_fu_39584_p3 = ((or_ln302_74_fu_39562_p2[0:0] == 1'b1) ? select_ln302_148_fu_39568_p3 : select_ln350_74_fu_39576_p3);

assign select_ln302_14_fu_23298_p3 = ((xor_ln302_14_fu_23280_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_255_fu_23242_p2);

assign select_ln302_150_fu_39670_p3 = ((xor_ln302_150_fu_39652_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_391_fu_39614_p2);

assign select_ln302_151_fu_39686_p3 = ((or_ln302_75_fu_39664_p2[0:0] == 1'b1) ? select_ln302_150_fu_39670_p3 : select_ln350_75_fu_39678_p3);

assign select_ln302_152_fu_39772_p3 = ((xor_ln302_152_fu_39754_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_393_fu_39716_p2);

assign select_ln302_153_fu_39788_p3 = ((or_ln302_76_fu_39766_p2[0:0] == 1'b1) ? select_ln302_152_fu_39772_p3 : select_ln350_76_fu_39780_p3);

assign select_ln302_154_fu_39874_p3 = ((xor_ln302_154_fu_39856_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_395_fu_39818_p2);

assign select_ln302_155_fu_39890_p3 = ((or_ln302_77_fu_39868_p2[0:0] == 1'b1) ? select_ln302_154_fu_39874_p3 : select_ln350_77_fu_39882_p3);

assign select_ln302_156_fu_39976_p3 = ((xor_ln302_156_fu_39958_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_397_fu_39920_p2);

assign select_ln302_157_fu_39992_p3 = ((or_ln302_78_fu_39970_p2[0:0] == 1'b1) ? select_ln302_156_fu_39976_p3 : select_ln350_78_fu_39984_p3);

assign select_ln302_158_fu_40078_p3 = ((xor_ln302_158_fu_40060_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_399_fu_40022_p2);

assign select_ln302_159_fu_40094_p3 = ((or_ln302_79_fu_40072_p2[0:0] == 1'b1) ? select_ln302_158_fu_40078_p3 : select_ln350_79_fu_40086_p3);

assign select_ln302_160_fu_40180_p3 = ((xor_ln302_160_fu_40162_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_401_fu_40124_p2);

assign select_ln302_161_fu_40196_p3 = ((or_ln302_80_fu_40174_p2[0:0] == 1'b1) ? select_ln302_160_fu_40180_p3 : select_ln350_80_fu_40188_p3);

assign select_ln302_16_fu_23396_p3 = ((xor_ln302_16_fu_23378_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_257_fu_23340_p2);

assign select_ln302_18_fu_23498_p3 = ((xor_ln302_18_fu_23480_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_259_fu_23442_p2);

assign select_ln302_20_fu_23600_p3 = ((xor_ln302_20_fu_23582_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_261_fu_23544_p2);

assign select_ln302_22_fu_23702_p3 = ((xor_ln302_22_fu_23684_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_263_fu_23646_p2);

assign select_ln302_24_fu_23804_p3 = ((xor_ln302_24_fu_23786_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_265_fu_23748_p2);

assign select_ln302_26_fu_23906_p3 = ((xor_ln302_26_fu_23888_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_267_fu_23850_p2);

assign select_ln302_28_fu_24008_p3 = ((xor_ln302_28_fu_23990_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_269_fu_23952_p2);

assign select_ln302_2_fu_22710_p3 = ((xor_ln302_2_fu_22692_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_243_fu_22654_p2);

assign select_ln302_30_fu_24110_p3 = ((xor_ln302_30_fu_24092_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_271_fu_24054_p2);

assign select_ln302_32_fu_24212_p3 = ((xor_ln302_32_fu_24194_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_273_fu_24156_p2);

assign select_ln302_34_fu_24314_p3 = ((xor_ln302_34_fu_24296_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_275_fu_24258_p2);

assign select_ln302_36_fu_28499_p3 = ((xor_ln302_36_fu_28481_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_277_fu_28444_p2);

assign select_ln302_38_fu_28599_p3 = ((xor_ln302_38_fu_28581_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_279_fu_28544_p2);

assign select_ln302_40_fu_28659_p3 = ((xor_ln302_40_fu_28643_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_281_reg_41723);

assign select_ln302_42_fu_28757_p3 = ((xor_ln302_42_fu_28739_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_283_fu_28702_p2);

assign select_ln302_44_fu_28857_p3 = ((xor_ln302_44_fu_28839_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_285_fu_28802_p2);

assign select_ln302_46_fu_28957_p3 = ((xor_ln302_46_fu_28939_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_287_fu_28902_p2);

assign select_ln302_48_fu_29017_p3 = ((xor_ln302_48_fu_29001_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_289_reg_41743);

assign select_ln302_4_fu_22808_p3 = ((xor_ln302_4_fu_22790_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_245_fu_22752_p2);

assign select_ln302_50_fu_29115_p3 = ((xor_ln302_50_fu_29097_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_291_fu_29060_p2);

assign select_ln302_52_fu_29215_p3 = ((xor_ln302_52_fu_29197_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_293_fu_29160_p2);

assign select_ln302_54_fu_29317_p3 = ((xor_ln302_54_fu_29299_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_295_fu_29261_p2);

assign select_ln302_56_fu_29419_p3 = ((xor_ln302_56_fu_29401_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_297_fu_29363_p2);

assign select_ln302_58_fu_29521_p3 = ((xor_ln302_58_fu_29503_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_299_fu_29465_p2);

assign select_ln302_60_fu_29623_p3 = ((xor_ln302_60_fu_29605_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_301_fu_29567_p2);

assign select_ln302_62_fu_29725_p3 = ((xor_ln302_62_fu_29707_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_303_fu_29669_p2);

assign select_ln302_64_fu_29827_p3 = ((xor_ln302_64_fu_29809_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_305_fu_29771_p2);

assign select_ln302_66_fu_29929_p3 = ((xor_ln302_66_fu_29911_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_307_fu_29873_p2);

assign select_ln302_68_fu_30031_p3 = ((xor_ln302_68_fu_30013_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_309_fu_29975_p2);

assign select_ln302_6_fu_22906_p3 = ((xor_ln302_6_fu_22888_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_247_fu_22850_p2);

assign select_ln302_70_fu_30133_p3 = ((xor_ln302_70_fu_30115_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_311_fu_30077_p2);

assign select_ln302_72_fu_33958_p3 = ((xor_ln302_72_fu_33942_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_313_reg_42241);

assign select_ln302_74_fu_34016_p3 = ((xor_ln302_74_fu_34000_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_315_reg_42261);

assign select_ln302_76_fu_30307_p3 = ((xor_ln302_76_fu_30289_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_317_fu_30251_p2);

assign select_ln302_78_fu_34074_p3 = ((xor_ln302_78_fu_34058_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_319_reg_42287);

assign select_ln302_80_fu_34132_p3 = ((xor_ln302_80_fu_34116_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_321_reg_42307);

assign select_ln302_82_fu_34190_p3 = ((xor_ln302_82_fu_34174_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_323_reg_42327);

assign select_ln302_84_fu_30517_p3 = ((xor_ln302_84_fu_30499_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_325_fu_30461_p2);

assign select_ln302_86_fu_34248_p3 = ((xor_ln302_86_fu_34232_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_327_reg_42353);

assign select_ln302_88_fu_34306_p3 = ((xor_ln302_88_fu_34290_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_329_reg_42373);

assign select_ln302_8_fu_23004_p3 = ((xor_ln302_8_fu_22986_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_249_fu_22948_p2);

assign select_ln302_90_fu_34406_p3 = ((xor_ln302_90_fu_34388_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_331_fu_34350_p2);

assign select_ln302_92_fu_34508_p3 = ((xor_ln302_92_fu_34490_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_333_fu_34452_p2);

assign select_ln302_94_fu_34608_p3 = ((xor_ln302_94_fu_34590_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_335_fu_34553_p2);

assign select_ln302_96_fu_34710_p3 = ((xor_ln302_96_fu_34692_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_337_fu_34654_p2);

assign select_ln302_98_fu_34812_p3 = ((xor_ln302_98_fu_34794_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_339_fu_34756_p2);

assign select_ln302_fu_22612_p3 = ((xor_ln302_fu_22594_p2[0:0] == 1'b1) ? 32'd2147483647 : p_Val2_241_fu_22556_p2);

assign select_ln346_100_fu_31233_p3 = ((overflow_50_fu_31204_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_102_fu_31258_p3 = ((overflow_51_reg_41931[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_104_fu_31375_p3 = ((overflow_52_fu_31346_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_106_fu_31400_p3 = ((overflow_53_reg_41977[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_108_fu_31541_p3 = ((overflow_54_fu_31512_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_10_fu_19109_p3 = ((overflow_5_fu_19080_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_110_fu_31690_p3 = ((overflow_55_fu_31661_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_112_fu_31839_p3 = ((overflow_56_fu_31810_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_114_fu_31988_p3 = ((overflow_57_fu_31959_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_116_fu_32137_p3 = ((overflow_58_fu_32108_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_118_fu_32286_p3 = ((overflow_59_fu_32257_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_120_fu_32435_p3 = ((overflow_60_fu_32406_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_122_fu_32460_p3 = ((overflow_61_reg_42195[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_124_fu_32601_p3 = ((overflow_62_fu_32572_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_126_fu_36263_p3 = ((overflow_63_fu_36234_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_128_fu_36388_p3 = ((overflow_64_fu_36359_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_12_fu_19134_p3 = ((overflow_6_reg_40498[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_130_fu_36513_p3 = ((overflow_65_fu_36484_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_132_fu_36638_p3 = ((overflow_66_fu_36609_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_134_fu_36763_p3 = ((overflow_67_fu_36734_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_136_fu_36788_p3 = ((overflow_68_reg_42546[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_138_fu_36905_p3 = ((overflow_69_fu_36876_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_140_fu_37030_p3 = ((overflow_70_fu_37001_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_142_fu_37155_p3 = ((overflow_71_fu_37126_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_144_fu_37304_p3 = ((overflow_72_fu_37275_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_146_fu_37453_p3 = ((overflow_73_fu_37424_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_148_fu_37602_p3 = ((overflow_74_fu_37573_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_14_fu_19248_p3 = ((overflow_7_fu_19219_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_150_fu_37751_p3 = ((overflow_75_fu_37722_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_152_fu_37776_p3 = ((overflow_76_reg_42770[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_154_fu_37917_p3 = ((overflow_77_fu_37888_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_156_fu_38066_p3 = ((overflow_78_fu_38037_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_158_fu_38215_p3 = ((overflow_79_fu_38186_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_160_fu_38364_p3 = ((overflow_80_fu_38335_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_16_fu_19372_p3 = ((overflow_8_fu_19343_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_18_fu_19521_p3 = ((overflow_9_fu_19492_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_20_fu_19546_p3 = ((overflow_10_reg_40604[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_22_fu_19563_p3 = ((overflow_11_reg_40619[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_24_fu_19704_p3 = ((overflow_12_fu_19675_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_26_fu_19853_p3 = ((overflow_13_fu_19824_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_28_fu_19878_p3 = ((overflow_14_reg_40692[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_2_fu_18717_p3 = ((overflow_1_fu_18688_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_30_fu_19995_p3 = ((overflow_15_fu_19966_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_32_fu_20144_p3 = ((overflow_16_fu_20115_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_34_fu_20293_p3 = ((overflow_17_fu_20264_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_36_fu_24413_p3 = ((overflow_18_reg_41048[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_38_fu_24430_p3 = ((overflow_19_reg_41063[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_40_fu_20700_p3 = ((overflow_20_fu_20671_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_42_fu_24447_p3 = ((overflow_21_reg_41078[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_44_fu_24464_p3 = ((overflow_22_reg_41093[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_46_fu_24481_p3 = ((overflow_23_reg_41108[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_48_fu_21112_p3 = ((overflow_24_reg_40970[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_4_fu_18742_p3 = ((overflow_2_reg_40390[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_50_fu_24498_p3 = ((overflow_25_reg_41123[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_52_fu_24515_p3 = ((overflow_26_reg_41138[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_54_fu_24629_p3 = ((overflow_27_fu_24600_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_56_fu_24753_p3 = ((overflow_28_fu_24724_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_58_fu_24878_p3 = ((overflow_29_fu_24849_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_60_fu_25003_p3 = ((overflow_30_fu_24974_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_62_fu_25128_p3 = ((overflow_31_fu_25099_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_64_fu_25253_p3 = ((overflow_32_fu_25224_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_66_fu_25378_p3 = ((overflow_33_fu_25349_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_68_fu_25503_p3 = ((overflow_34_fu_25474_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_6_fu_18859_p3 = ((overflow_3_fu_18830_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_70_fu_25625_p3 = ((overflow_35_fu_25596_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_72_fu_25773_p3 = ((overflow_36_fu_25744_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_74_fu_25922_p3 = ((overflow_37_fu_25893_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_76_fu_26071_p3 = ((overflow_38_fu_26042_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_78_fu_26096_p3 = ((overflow_39_reg_41519[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_80_fu_26237_p3 = ((overflow_40_fu_26208_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_82_fu_26386_p3 = ((overflow_41_fu_26357_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_84_fu_26535_p3 = ((overflow_42_fu_26506_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_86_fu_26684_p3 = ((overflow_43_fu_26655_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_88_fu_26833_p3 = ((overflow_44_fu_26804_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_8_fu_18984_p3 = ((overflow_4_fu_18955_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_90_fu_30616_p3 = ((overflow_45_reg_41761[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_92_fu_30733_p3 = ((overflow_46_fu_30704_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_94_fu_30858_p3 = ((overflow_47_fu_30829_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_96_fu_30983_p3 = ((overflow_48_fu_30954_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_98_fu_31108_p3 = ((overflow_49_fu_31079_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln346_fu_18592_p3 = ((overflow_fu_18563_p2[0:0] == 1'b1) ? 32'd2147483647 : 32'd2147483648);

assign select_ln350_10_fu_23608_p3 = ((underflow_91_fu_23576_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_261_fu_23544_p2);

assign select_ln350_11_fu_23710_p3 = ((underflow_92_fu_23678_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_263_fu_23646_p2);

assign select_ln350_12_fu_23812_p3 = ((underflow_93_fu_23780_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_265_fu_23748_p2);

assign select_ln350_13_fu_23914_p3 = ((underflow_94_fu_23882_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_267_fu_23850_p2);

assign select_ln350_14_fu_24016_p3 = ((underflow_95_fu_23984_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_269_fu_23952_p2);

assign select_ln350_15_fu_24118_p3 = ((underflow_96_fu_24086_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_271_fu_24054_p2);

assign select_ln350_16_fu_24220_p3 = ((underflow_97_fu_24188_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_273_fu_24156_p2);

assign select_ln350_17_fu_24322_p3 = ((underflow_98_fu_24290_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_275_fu_24258_p2);

assign select_ln350_18_fu_28507_p3 = ((underflow_99_fu_28475_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_277_fu_28444_p2);

assign select_ln350_19_fu_28607_p3 = ((underflow_100_fu_28575_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_279_fu_28544_p2);

assign select_ln350_1_fu_22718_p3 = ((underflow_82_fu_22686_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_243_fu_22654_p2);

assign select_ln350_20_fu_28666_p3 = ((underflow_101_fu_28638_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_281_reg_41723);

assign select_ln350_21_fu_28765_p3 = ((underflow_102_fu_28733_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_283_fu_28702_p2);

assign select_ln350_22_fu_28865_p3 = ((underflow_103_fu_28833_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_285_fu_28802_p2);

assign select_ln350_23_fu_28965_p3 = ((underflow_104_fu_28933_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_287_fu_28902_p2);

assign select_ln350_24_fu_29024_p3 = ((underflow_105_fu_28996_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_289_reg_41743);

assign select_ln350_25_fu_29123_p3 = ((underflow_106_fu_29091_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_291_fu_29060_p2);

assign select_ln350_26_fu_29223_p3 = ((underflow_107_fu_29191_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_293_fu_29160_p2);

assign select_ln350_27_fu_29325_p3 = ((underflow_108_fu_29293_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_295_fu_29261_p2);

assign select_ln350_28_fu_29427_p3 = ((underflow_109_fu_29395_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_297_fu_29363_p2);

assign select_ln350_29_fu_29529_p3 = ((underflow_110_fu_29497_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_299_fu_29465_p2);

assign select_ln350_2_fu_22816_p3 = ((underflow_83_fu_22784_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_245_fu_22752_p2);

assign select_ln350_30_fu_29631_p3 = ((underflow_111_fu_29599_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_301_fu_29567_p2);

assign select_ln350_31_fu_29733_p3 = ((underflow_112_fu_29701_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_303_fu_29669_p2);

assign select_ln350_32_fu_29835_p3 = ((underflow_113_fu_29803_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_305_fu_29771_p2);

assign select_ln350_33_fu_29937_p3 = ((underflow_114_fu_29905_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_307_fu_29873_p2);

assign select_ln350_34_fu_30039_p3 = ((underflow_115_fu_30007_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_309_fu_29975_p2);

assign select_ln350_35_fu_30141_p3 = ((underflow_116_fu_30109_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_311_fu_30077_p2);

assign select_ln350_36_fu_33965_p3 = ((underflow_117_fu_33937_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_313_reg_42241);

assign select_ln350_37_fu_34023_p3 = ((underflow_118_fu_33995_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_315_reg_42261);

assign select_ln350_38_fu_30315_p3 = ((underflow_119_fu_30283_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_317_fu_30251_p2);

assign select_ln350_39_fu_34081_p3 = ((underflow_120_fu_34053_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_319_reg_42287);

assign select_ln350_3_fu_22914_p3 = ((underflow_84_fu_22882_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_247_fu_22850_p2);

assign select_ln350_40_fu_34139_p3 = ((underflow_121_fu_34111_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_321_reg_42307);

assign select_ln350_41_fu_34197_p3 = ((underflow_122_fu_34169_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_323_reg_42327);

assign select_ln350_42_fu_30525_p3 = ((underflow_123_fu_30493_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_325_fu_30461_p2);

assign select_ln350_43_fu_34255_p3 = ((underflow_124_fu_34227_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_327_reg_42353);

assign select_ln350_44_fu_34313_p3 = ((underflow_125_fu_34285_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_329_reg_42373);

assign select_ln350_45_fu_34414_p3 = ((underflow_126_fu_34382_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_331_fu_34350_p2);

assign select_ln350_46_fu_34516_p3 = ((underflow_127_fu_34484_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_333_fu_34452_p2);

assign select_ln350_47_fu_34616_p3 = ((underflow_128_fu_34584_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_335_fu_34553_p2);

assign select_ln350_48_fu_34718_p3 = ((underflow_129_fu_34686_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_337_fu_34654_p2);

assign select_ln350_49_fu_34820_p3 = ((underflow_130_fu_34788_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_339_fu_34756_p2);

assign select_ln350_4_fu_23012_p3 = ((underflow_85_fu_22980_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_249_fu_22948_p2);

assign select_ln350_50_fu_34922_p3 = ((underflow_131_fu_34890_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_341_fu_34858_p2);

assign select_ln350_51_fu_35022_p3 = ((underflow_132_fu_34990_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_343_fu_34959_p2);

assign select_ln350_52_fu_35124_p3 = ((underflow_133_fu_35092_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_345_fu_35060_p2);

assign select_ln350_53_fu_35226_p3 = ((underflow_134_fu_35194_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_347_fu_35162_p2);

assign select_ln350_54_fu_35328_p3 = ((underflow_135_fu_35296_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_349_fu_35264_p2);

assign select_ln350_55_fu_35430_p3 = ((underflow_136_fu_35398_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_351_fu_35366_p2);

assign select_ln350_56_fu_35532_p3 = ((underflow_137_fu_35500_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_353_fu_35468_p2);

assign select_ln350_57_fu_35634_p3 = ((underflow_138_fu_35602_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_355_fu_35570_p2);

assign select_ln350_58_fu_35736_p3 = ((underflow_139_fu_35704_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_357_fu_35672_p2);

assign select_ln350_59_fu_35838_p3 = ((underflow_140_fu_35806_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_359_fu_35774_p2);

assign select_ln350_5_fu_23110_p3 = ((underflow_86_fu_23078_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_251_fu_23046_p2);

assign select_ln350_60_fu_35940_p3 = ((underflow_141_fu_35908_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_361_fu_35876_p2);

assign select_ln350_61_fu_36042_p3 = ((underflow_142_fu_36010_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_363_fu_35978_p2);

assign select_ln350_62_fu_36144_p3 = ((underflow_143_fu_36112_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_365_fu_36080_p2);

assign select_ln350_63_fu_38470_p3 = ((underflow_144_fu_38438_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_367_fu_38407_p2);

assign select_ln350_64_fu_38570_p3 = ((underflow_145_fu_38538_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_369_fu_38507_p2);

assign select_ln350_65_fu_38670_p3 = ((underflow_146_fu_38638_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_371_fu_38607_p2);

assign select_ln350_66_fu_38770_p3 = ((underflow_147_fu_38738_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_373_fu_38707_p2);

assign select_ln350_67_fu_38870_p3 = ((underflow_148_fu_38838_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_375_fu_38807_p2);

assign select_ln350_68_fu_38970_p3 = ((underflow_149_fu_38938_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_377_fu_38907_p2);

assign select_ln350_69_fu_39070_p3 = ((underflow_150_fu_39038_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_379_fu_39007_p2);

assign select_ln350_6_fu_23208_p3 = ((underflow_87_fu_23176_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_253_fu_23144_p2);

assign select_ln350_70_fu_39170_p3 = ((underflow_151_fu_39138_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_381_fu_39107_p2);

assign select_ln350_71_fu_39270_p3 = ((underflow_152_fu_39238_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_383_fu_39207_p2);

assign select_ln350_72_fu_39372_p3 = ((underflow_153_fu_39340_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_385_fu_39308_p2);

assign select_ln350_73_fu_39474_p3 = ((underflow_154_fu_39442_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_387_fu_39410_p2);

assign select_ln350_74_fu_39576_p3 = ((underflow_155_fu_39544_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_389_fu_39512_p2);

assign select_ln350_75_fu_39678_p3 = ((underflow_156_fu_39646_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_391_fu_39614_p2);

assign select_ln350_76_fu_39780_p3 = ((underflow_157_fu_39748_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_393_fu_39716_p2);

assign select_ln350_77_fu_39882_p3 = ((underflow_158_fu_39850_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_395_fu_39818_p2);

assign select_ln350_78_fu_39984_p3 = ((underflow_159_fu_39952_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_397_fu_39920_p2);

assign select_ln350_79_fu_40086_p3 = ((underflow_160_fu_40054_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_399_fu_40022_p2);

assign select_ln350_7_fu_23306_p3 = ((underflow_88_fu_23274_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_255_fu_23242_p2);

assign select_ln350_80_fu_40188_p3 = ((underflow_161_fu_40156_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_401_fu_40124_p2);

assign select_ln350_8_fu_23404_p3 = ((underflow_89_fu_23372_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_257_fu_23340_p2);

assign select_ln350_9_fu_23506_p3 = ((underflow_90_fu_23474_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_259_fu_23442_p2);

assign select_ln350_fu_22620_p3 = ((underflow_81_fu_22588_p2[0:0] == 1'b1) ? 32'd2147483648 : p_Val2_241_fu_22556_p2);

assign sext_ln1273_10_fu_32967_p1 = $signed(shl_ln1273_s_fu_32960_p3);

assign sext_ln1273_11_fu_33553_p1 = $signed(shl_ln1273_10_fu_33546_p3);

assign sext_ln1273_12_fu_33564_p1 = $signed(shl_ln1273_11_fu_33557_p3);

assign sext_ln1273_1_fu_18177_p1 = $signed(shl_ln1273_1_fu_18169_p3);

assign sext_ln1273_2_fu_18189_p1 = $signed(shl_ln1273_2_fu_18181_p3);

assign sext_ln1273_3_fu_22138_p1 = $signed(shl_ln1273_3_fu_22131_p3);

assign sext_ln1273_4_fu_26883_p1 = $signed(shl_ln1273_4_fu_26876_p3);

assign sext_ln1273_5_fu_27391_p1 = $signed(shl_ln1273_5_fu_27384_p3);

assign sext_ln1273_6_fu_27408_p1 = $signed(shl_ln1273_6_fu_27401_p3);

assign sext_ln1273_7_fu_27669_p1 = $signed(shl_ln1273_7_fu_27662_p3);

assign sext_ln1273_8_fu_28180_p1 = $signed(shl_ln1273_8_fu_28173_p3);

assign sext_ln1273_9_fu_28191_p1 = $signed(shl_ln1273_9_fu_28184_p3);

assign sext_ln1273_fu_16419_p1 = $signed(shl_ln_fu_16411_p3);

assign sext_ln70_13_fu_17909_p0 = p_read2_int_reg;

assign sext_ln70_13_fu_17909_p1 = sext_ln70_13_fu_17909_p0;

assign sext_ln70_15_fu_21388_p1 = p_read_23_reg_40314;

assign sext_ln70_16_fu_21393_p1 = p_read_23_reg_40314;

assign sext_ln70_17_fu_21398_p1 = p_read_23_reg_40314;

assign sext_ln70_18_fu_21403_p1 = p_read_23_reg_40314;

assign sext_ln70_1_fu_16257_p0 = p_read_int_reg;

assign sext_ln70_1_fu_16257_p1 = sext_ln70_1_fu_16257_p0;

assign sext_ln70_21_fu_21984_p1 = p_read_22_reg_40302;

assign sext_ln70_22_fu_21989_p1 = p_read_22_reg_40302;

assign sext_ln70_24_fu_21996_p1 = p_read_22_reg_40302;

assign sext_ln70_29_fu_26867_p1 = p_read_21_reg_40289_pp0_iter1_reg;

assign sext_ln70_2_fu_16263_p0 = p_read_int_reg;

assign sext_ln70_2_fu_16263_p1 = sext_ln70_2_fu_16263_p0;

assign sext_ln70_30_fu_26873_p1 = p_read_21_reg_40289_pp0_iter1_reg;

assign sext_ln70_31_fu_27859_p1 = p_read_20_reg_40279_pp0_iter1_reg;

assign sext_ln70_32_fu_27865_p1 = p_read_20_reg_40279_pp0_iter1_reg;

assign sext_ln70_35_fu_32623_p1 = p_read_19_reg_40271_pp0_iter2_reg;

assign sext_ln70_36_fu_32629_p1 = p_read_19_reg_40271_pp0_iter2_reg;

assign sext_ln70_37_fu_32634_p1 = p_read_19_reg_40271_pp0_iter2_reg;

assign sext_ln70_3_fu_16269_p0 = p_read_int_reg;

assign sext_ln70_3_fu_16269_p1 = sext_ln70_3_fu_16269_p0;

assign sext_ln70_43_fu_33369_p1 = p_read_18_reg_40258_pp0_iter2_reg;

assign sext_ln70_7_fu_17134_p0 = p_read1_int_reg;

assign sext_ln70_7_fu_17134_p1 = sext_ln70_7_fu_17134_p0;

assign sext_ln70_8_fu_17141_p0 = p_read1_int_reg;

assign sext_ln70_8_fu_17141_p1 = sext_ln70_8_fu_17141_p0;

assign sext_ln813_100_fu_35246_p1 = rhs_54_fu_31555_p3;

assign sext_ln813_101_fu_35344_p1 = lhs_46_fu_34524_p3;

assign sext_ln813_102_fu_35348_p1 = rhs_55_fu_31704_p3;

assign sext_ln813_103_fu_35446_p1 = lhs_47_fu_34624_p3;

assign sext_ln813_104_fu_35450_p1 = rhs_56_fu_31853_p3;

assign sext_ln813_105_fu_35548_p1 = lhs_48_fu_34726_p3;

assign sext_ln813_106_fu_35552_p1 = rhs_57_fu_32002_p3;

assign sext_ln813_107_fu_35650_p1 = lhs_49_fu_34828_p3;

assign sext_ln813_108_fu_35654_p1 = rhs_58_fu_32151_p3;

assign sext_ln813_109_fu_35752_p1 = lhs_50_fu_34930_p3;

assign sext_ln813_10_fu_23424_p1 = rhs_9_fu_19535_p3;

assign sext_ln813_110_fu_35756_p1 = rhs_59_fu_32300_p3;

assign sext_ln813_111_fu_35854_p1 = lhs_51_fu_35030_p3;

assign sext_ln813_112_fu_35858_p1 = rhs_60_fu_32449_p3;

assign sext_ln813_113_fu_35956_p1 = lhs_52_fu_35132_p3;

assign sext_ln813_114_fu_35960_p1 = rhs_61_fu_32467_p3;

assign sext_ln813_115_fu_36058_p1 = lhs_53_fu_35234_p3;

assign sext_ln813_116_fu_36062_p1 = rhs_62_fu_32615_p3;

assign sext_ln813_117_fu_38386_p1 = lhs_54_reg_42896;

assign sext_ln813_118_fu_38389_p1 = rhs_63_fu_36277_p3;

assign sext_ln813_119_fu_38486_p1 = lhs_55_reg_42902;

assign sext_ln813_11_fu_23522_p1 = lhs_1_fu_22726_p3;

assign sext_ln813_120_fu_38489_p1 = rhs_64_fu_36402_p3;

assign sext_ln813_121_fu_38586_p1 = lhs_56_reg_42908;

assign sext_ln813_122_fu_38589_p1 = rhs_65_fu_36527_p3;

assign sext_ln813_123_fu_38686_p1 = lhs_57_reg_42914;

assign sext_ln813_124_fu_38689_p1 = rhs_66_fu_36652_p3;

assign sext_ln813_125_fu_38786_p1 = lhs_58_reg_42920;

assign sext_ln813_126_fu_38789_p1 = rhs_67_fu_36777_p3;

assign sext_ln813_127_fu_38886_p1 = lhs_59_reg_42926;

assign sext_ln813_128_fu_38889_p1 = rhs_68_fu_36795_p3;

assign sext_ln813_129_fu_38986_p1 = lhs_60_reg_42932;

assign sext_ln813_12_fu_23526_p1 = rhs_10_fu_19553_p3;

assign sext_ln813_130_fu_38989_p1 = rhs_69_fu_36919_p3;

assign sext_ln813_131_fu_39086_p1 = lhs_61_reg_42938;

assign sext_ln813_132_fu_39089_p1 = rhs_70_fu_37044_p3;

assign sext_ln813_133_fu_39186_p1 = lhs_62_reg_42944;

assign sext_ln813_134_fu_39189_p1 = rhs_71_fu_37169_p3;

assign sext_ln813_135_fu_39286_p1 = lhs_63_fu_38478_p3;

assign sext_ln813_136_fu_39290_p1 = rhs_72_fu_37318_p3;

assign sext_ln813_137_fu_39388_p1 = lhs_64_fu_38578_p3;

assign sext_ln813_138_fu_39392_p1 = rhs_73_fu_37467_p3;

assign sext_ln813_139_fu_39490_p1 = lhs_65_fu_38678_p3;

assign sext_ln813_13_fu_23624_p1 = lhs_2_fu_22824_p3;

assign sext_ln813_140_fu_39494_p1 = rhs_74_fu_37616_p3;

assign sext_ln813_141_fu_39592_p1 = lhs_66_fu_38778_p3;

assign sext_ln813_142_fu_39596_p1 = rhs_75_fu_37765_p3;

assign sext_ln813_143_fu_39694_p1 = lhs_67_fu_38878_p3;

assign sext_ln813_144_fu_39698_p1 = rhs_76_fu_37783_p3;

assign sext_ln813_145_fu_39796_p1 = lhs_68_fu_38978_p3;

assign sext_ln813_146_fu_39800_p1 = rhs_77_fu_37931_p3;

assign sext_ln813_147_fu_39898_p1 = lhs_69_fu_39078_p3;

assign sext_ln813_148_fu_39902_p1 = rhs_78_fu_38080_p3;

assign sext_ln813_149_fu_40000_p1 = lhs_70_fu_39178_p3;

assign sext_ln813_14_fu_23628_p1 = rhs_11_fu_19570_p3;

assign sext_ln813_150_fu_40004_p1 = rhs_79_fu_38229_p3;

assign sext_ln813_151_fu_40102_p1 = lhs_71_fu_39278_p3;

assign sext_ln813_152_fu_40106_p1 = rhs_80_fu_38378_p3;

assign sext_ln813_15_fu_23726_p1 = lhs_3_fu_22922_p3;

assign sext_ln813_16_fu_23730_p1 = rhs_12_fu_19718_p3;

assign sext_ln813_17_fu_23828_p1 = lhs_4_fu_23020_p3;

assign sext_ln813_18_fu_23832_p1 = rhs_13_fu_19867_p3;

assign sext_ln813_19_fu_23930_p1 = lhs_5_fu_23118_p3;

assign sext_ln813_1_fu_22636_p1 = rhs_1_fu_18731_p3;

assign sext_ln813_20_fu_23934_p1 = rhs_14_fu_19885_p3;

assign sext_ln813_21_fu_24032_p1 = lhs_6_fu_23216_p3;

assign sext_ln813_22_fu_24036_p1 = rhs_15_fu_20009_p3;

assign sext_ln813_23_fu_24134_p1 = lhs_7_fu_23314_p3;

assign sext_ln813_24_fu_24138_p1 = rhs_16_fu_20158_p3;

assign sext_ln813_25_fu_24236_p1 = lhs_8_fu_23412_p3;

assign sext_ln813_26_fu_24240_p1 = rhs_17_fu_20307_p3;

assign sext_ln813_27_fu_28423_p1 = lhs_9_reg_41674;

assign sext_ln813_28_fu_28426_p1 = rhs_18_fu_24420_p3;

assign sext_ln813_29_fu_28523_p1 = lhs_10_reg_41680;

assign sext_ln813_2_fu_22734_p1 = rhs_2_fu_18749_p3;

assign sext_ln813_30_fu_28526_p1 = rhs_19_fu_24437_p3;

assign sext_ln813_31_fu_24338_p1 = lhs_11_fu_23718_p3;

assign sext_ln813_32_fu_24342_p1 = rhs_20_fu_20714_p3;

assign sext_ln813_33_fu_28681_p1 = lhs_12_reg_41686;

assign sext_ln813_34_fu_28684_p1 = rhs_21_fu_24454_p3;

assign sext_ln813_35_fu_28781_p1 = lhs_13_reg_41692;

assign sext_ln813_36_fu_28784_p1 = rhs_22_fu_24471_p3;

assign sext_ln813_37_fu_28881_p1 = lhs_14_reg_41698;

assign sext_ln813_38_fu_28884_p1 = rhs_23_fu_24488_p3;

assign sext_ln813_39_fu_24374_p1 = lhs_15_fu_24126_p3;

assign sext_ln813_3_fu_22832_p1 = rhs_3_fu_18873_p3;

assign sext_ln813_40_fu_24378_p1 = rhs_24_fu_21119_p3;

assign sext_ln813_41_fu_29039_p1 = lhs_16_reg_41704;

assign sext_ln813_42_fu_29042_p1 = rhs_25_fu_24505_p3;

assign sext_ln813_43_fu_29139_p1 = lhs_17_reg_41710;

assign sext_ln813_44_fu_29142_p1 = rhs_26_fu_24522_p3;

assign sext_ln813_45_fu_29239_p1 = lhs_18_fu_28515_p3;

assign sext_ln813_46_fu_29243_p1 = rhs_27_fu_24643_p3;

assign sext_ln813_47_fu_29341_p1 = lhs_19_fu_28615_p3;

assign sext_ln813_48_fu_29345_p1 = rhs_28_fu_24767_p3;

assign sext_ln813_49_fu_29443_p1 = lhs_20_fu_28673_p3;

assign sext_ln813_4_fu_22930_p1 = rhs_4_fu_18998_p3;

assign sext_ln813_50_fu_29447_p1 = rhs_29_fu_24892_p3;

assign sext_ln813_51_fu_29545_p1 = lhs_21_fu_28773_p3;

assign sext_ln813_52_fu_29549_p1 = rhs_30_fu_25017_p3;

assign sext_ln813_53_fu_29647_p1 = lhs_22_fu_28873_p3;

assign sext_ln813_54_fu_29651_p1 = rhs_31_fu_25142_p3;

assign sext_ln813_55_fu_29749_p1 = lhs_23_fu_28973_p3;

assign sext_ln813_56_fu_29753_p1 = rhs_32_fu_25267_p3;

assign sext_ln813_57_fu_29851_p1 = lhs_24_fu_29031_p3;

assign sext_ln813_58_fu_29855_p1 = rhs_33_fu_25392_p3;

assign sext_ln813_59_fu_29953_p1 = lhs_25_fu_29131_p3;

assign sext_ln813_5_fu_23028_p1 = rhs_5_fu_19123_p3;

assign sext_ln813_60_fu_29957_p1 = rhs_34_fu_25517_p3;

assign sext_ln813_61_fu_30055_p1 = lhs_26_fu_29231_p3;

assign sext_ln813_62_fu_30059_p1 = rhs_35_fu_25639_p3;

assign sext_ln813_63_fu_30157_p1 = lhs_27_fu_29333_p3;

assign sext_ln813_64_fu_30161_p1 = rhs_36_fu_25787_p3;

assign sext_ln813_65_fu_30193_p1 = lhs_28_fu_29435_p3;

assign sext_ln813_66_fu_30197_p1 = rhs_37_fu_25936_p3;

assign sext_ln813_67_fu_30229_p1 = lhs_29_fu_29537_p3;

assign sext_ln813_68_fu_30233_p1 = rhs_38_fu_26085_p3;

assign sext_ln813_69_fu_30331_p1 = lhs_30_fu_29639_p3;

assign sext_ln813_6_fu_23126_p1 = rhs_6_fu_19141_p3;

assign sext_ln813_70_fu_30335_p1 = rhs_39_fu_26103_p3;

assign sext_ln813_71_fu_30367_p1 = lhs_31_fu_29741_p3;

assign sext_ln813_72_fu_30371_p1 = rhs_40_fu_26251_p3;

assign sext_ln813_73_fu_30403_p1 = lhs_32_fu_29843_p3;

assign sext_ln813_74_fu_30407_p1 = rhs_41_fu_26400_p3;

assign sext_ln813_75_fu_30439_p1 = lhs_33_fu_29945_p3;

assign sext_ln813_76_fu_30443_p1 = rhs_42_fu_26549_p3;

assign sext_ln813_77_fu_30541_p1 = lhs_34_fu_30047_p3;

assign sext_ln813_78_fu_30545_p1 = rhs_43_fu_26698_p3;

assign sext_ln813_79_fu_30577_p1 = lhs_35_fu_30149_p3;

assign sext_ln813_7_fu_23224_p1 = rhs_7_fu_19262_p3;

assign sext_ln813_80_fu_30581_p1 = rhs_44_fu_26847_p3;

assign sext_ln813_81_fu_34328_p1 = lhs_36_fu_33972_p3;

assign sext_ln813_82_fu_34332_p1 = rhs_45_fu_30623_p3;

assign sext_ln813_83_fu_34430_p1 = lhs_37_fu_34030_p3;

assign sext_ln813_84_fu_34434_p1 = rhs_46_fu_30747_p3;

assign sext_ln813_85_fu_34532_p1 = lhs_38_reg_42274;

assign sext_ln813_86_fu_34535_p1 = rhs_47_fu_30872_p3;

assign sext_ln813_87_fu_34632_p1 = lhs_39_fu_34088_p3;

assign sext_ln813_88_fu_34636_p1 = rhs_48_fu_30997_p3;

assign sext_ln813_89_fu_34734_p1 = lhs_40_fu_34146_p3;

assign sext_ln813_8_fu_23322_p1 = rhs_8_fu_19386_p3;

assign sext_ln813_90_fu_34738_p1 = rhs_49_fu_31122_p3;

assign sext_ln813_91_fu_34836_p1 = lhs_41_fu_34204_p3;

assign sext_ln813_92_fu_34840_p1 = rhs_50_fu_31247_p3;

assign sext_ln813_93_fu_34938_p1 = lhs_42_reg_42340;

assign sext_ln813_94_fu_34941_p1 = rhs_51_fu_31265_p3;

assign sext_ln813_95_fu_35038_p1 = lhs_43_fu_34262_p3;

assign sext_ln813_96_fu_35042_p1 = rhs_52_fu_31389_p3;

assign sext_ln813_97_fu_35140_p1 = lhs_44_fu_34320_p3;

assign sext_ln813_98_fu_35144_p1 = rhs_53_fu_31407_p3;

assign sext_ln813_99_fu_35242_p1 = lhs_45_fu_34422_p3;

assign sext_ln813_9_fu_23420_p1 = lhs_fu_22628_p3;

assign sext_ln813_fu_22538_p1 = rhs_fu_18606_p3;

assign sext_ln823_10_fu_17083_p1 = $signed(p_Val2_25_fu_17073_p4);

assign sext_ln823_11_fu_19394_p1 = $signed(p_Val2_28_reg_40576);

assign sext_ln823_12_fu_19577_p1 = $signed(p_Val2_35_reg_40635);

assign sext_ln823_13_fu_19726_p1 = $signed(p_Val2_38_reg_40664);

assign sext_ln823_14_fu_17759_p1 = $signed(p_Val2_43_fu_17749_p4);

assign sext_ln823_15_fu_20017_p1 = $signed(p_Val2_46_reg_40739);

assign sext_ln823_16_fu_20166_p1 = $signed(p_Val2_49_reg_40768);

assign sext_ln823_17_fu_20315_p1 = $signed(p_Val2_52_reg_40797);

assign sext_ln823_18_fu_20444_p1 = $signed(p_Val2_55_reg_40826);

assign sext_ln823_19_fu_20573_p1 = $signed(p_Val2_58_reg_40855);

assign sext_ln823_1_fu_17379_p1 = $signed(p_Val2_32_fu_17369_p4);

assign sext_ln823_20_fu_20722_p1 = $signed(p_Val2_61_reg_40884);

assign sext_ln823_21_fu_20851_p1 = $signed(p_Val2_64_reg_40913);

assign sext_ln823_22_fu_20980_p1 = $signed(p_Val2_67_reg_40942);

assign sext_ln823_23_fu_18217_p1 = $signed(p_Val2_70_fu_18207_p4);

assign sext_ln823_24_fu_21126_p1 = $signed(p_Val2_73_reg_40986);

assign sext_ln823_25_fu_21255_p1 = $signed(p_Val2_76_reg_41015);

assign sext_ln823_26_fu_21486_p1 = $signed(p_Val2_82_fu_21476_p4);

assign sext_ln823_27_fu_21550_p1 = $signed(p_Val2_85_fu_21540_p4);

assign sext_ln823_28_fu_21614_p1 = $signed(p_Val2_88_fu_21604_p4);

assign sext_ln823_29_fu_21678_p1 = $signed(p_Val2_91_fu_21668_p4);

assign sext_ln823_2_fu_17607_p1 = $signed(p_Val2_40_fu_17597_p4);

assign sext_ln823_30_fu_21742_p1 = $signed(p_Val2_94_fu_21732_p4);

assign sext_ln823_31_fu_21806_p1 = $signed(p_Val2_97_fu_21796_p4);

assign sext_ln823_32_fu_21870_p1 = $signed(p_Val2_100_fu_21860_p4);

assign sext_ln823_33_fu_25646_p1 = $signed(p_Val2_106_reg_41433);

assign sext_ln823_34_fu_25795_p1 = $signed(p_Val2_109_reg_41462);

assign sext_ln823_35_fu_25944_p1 = $signed(p_Val2_112_reg_41491);

assign sext_ln823_36_fu_22166_p1 = $signed(p_Val2_115_fu_22156_p4);

assign sext_ln823_37_fu_26110_p1 = $signed(p_Val2_118_reg_41535);

assign sext_ln823_38_fu_26259_p1 = $signed(p_Val2_121_reg_41564);

assign sext_ln823_39_fu_26408_p1 = $signed(p_Val2_124_reg_41593);

assign sext_ln823_3_fu_16301_p1 = $signed(p_Val2_1_fu_16291_p4);

assign sext_ln823_40_fu_26557_p1 = $signed(p_Val2_127_reg_41622);

assign sext_ln823_41_fu_26706_p1 = $signed(p_Val2_130_reg_41651);

assign sext_ln823_42_fu_26911_p1 = $signed(p_Val2_133_fu_26901_p4);

assign sext_ln823_43_fu_27082_p1 = $signed(p_Val2_136_fu_27072_p4);

assign sext_ln823_44_fu_27146_p1 = $signed(p_Val2_139_fu_27136_p4);

assign sext_ln823_45_fu_27210_p1 = $signed(p_Val2_142_fu_27200_p4);

assign sext_ln823_46_fu_27274_p1 = $signed(p_Val2_145_fu_27264_p4);

assign sext_ln823_47_fu_27338_p1 = $signed(p_Val2_148_fu_27328_p4);

assign sext_ln823_48_fu_27436_p1 = $signed(p_Val2_151_fu_27426_p4);

assign sext_ln823_49_fu_27616_p1 = $signed(p_Val2_154_fu_27606_p4);

assign sext_ln823_4_fu_16365_p1 = $signed(p_Val2_4_fu_16355_p4);

assign sext_ln823_50_fu_27697_p1 = $signed(p_Val2_157_fu_27687_p4);

assign sext_ln823_51_fu_31414_p1 = $signed(p_Val2_160_reg_41993);

assign sext_ln823_52_fu_31563_p1 = $signed(p_Val2_163_reg_42022);

assign sext_ln823_53_fu_31712_p1 = $signed(p_Val2_166_reg_42051);

assign sext_ln823_54_fu_31861_p1 = $signed(p_Val2_169_reg_42080);

assign sext_ln823_55_fu_32010_p1 = $signed(p_Val2_172_reg_42109);

assign sext_ln823_56_fu_32159_p1 = $signed(p_Val2_175_reg_42138);

assign sext_ln823_57_fu_32308_p1 = $signed(p_Val2_178_reg_42167);

assign sext_ln823_58_fu_28219_p1 = $signed(p_Val2_181_fu_28209_p4);

assign sext_ln823_59_fu_32474_p1 = $signed(p_Val2_184_reg_42211);

assign sext_ln823_5_fu_16459_p1 = $signed(p_Val2_7_fu_16449_p4);

assign sext_ln823_60_fu_32658_p1 = $signed(p_Val2_187_fu_32648_p4);

assign sext_ln823_61_fu_32722_p1 = $signed(p_Val2_190_fu_32712_p4);

assign sext_ln823_62_fu_32786_p1 = $signed(p_Val2_193_fu_32776_p4);

assign sext_ln823_63_fu_32850_p1 = $signed(p_Val2_196_fu_32840_p4);

assign sext_ln823_64_fu_32914_p1 = $signed(p_Val2_199_fu_32904_p4);

assign sext_ln823_65_fu_32995_p1 = $signed(p_Val2_202_fu_32985_p4);

assign sext_ln823_66_fu_33175_p1 = $signed(p_Val2_205_fu_33165_p4);

assign sext_ln823_67_fu_33239_p1 = $signed(p_Val2_208_fu_33229_p4);

assign sext_ln823_68_fu_33303_p1 = $signed(p_Val2_211_fu_33293_p4);

assign sext_ln823_69_fu_37177_p1 = $signed(p_Val2_214_reg_42655);

assign sext_ln823_6_fu_16645_p1 = $signed(p_Val2_10_fu_16635_p4);

assign sext_ln823_70_fu_37326_p1 = $signed(p_Val2_217_reg_42684);

assign sext_ln823_71_fu_37475_p1 = $signed(p_Val2_220_reg_42713);

assign sext_ln823_72_fu_37624_p1 = $signed(p_Val2_223_reg_42742);

assign sext_ln823_73_fu_33592_p1 = $signed(p_Val2_226_fu_33582_p4);

assign sext_ln823_74_fu_37790_p1 = $signed(p_Val2_229_reg_42786);

assign sext_ln823_75_fu_37939_p1 = $signed(p_Val2_232_reg_42815);

assign sext_ln823_76_fu_38088_p1 = $signed(p_Val2_235_reg_42844);

assign sext_ln823_77_fu_38237_p1 = $signed(p_Val2_238_reg_42873);

assign sext_ln823_7_fu_16709_p1 = $signed(p_Val2_13_fu_16699_p4);

assign sext_ln823_8_fu_16773_p1 = $signed(p_Val2_16_fu_16763_p4);

assign sext_ln823_9_fu_16843_p1 = $signed(p_Val2_19_fu_16833_p4);

assign sext_ln823_fu_17207_p1 = $signed(p_Val2_30_fu_17197_p4);

assign sext_ln856_10_fu_19269_p1 = p_Val2_26_reg_40551;

assign sext_ln856_11_fu_19406_p1 = p_Val2_29_fu_19400_p2;

assign sext_ln856_12_fu_19589_p1 = p_Val2_36_fu_19583_p2;

assign sext_ln856_13_fu_19738_p1 = p_Val2_39_fu_19732_p2;

assign sext_ln856_14_fu_19892_p1 = p_Val2_44_reg_40714;

assign sext_ln856_15_fu_20029_p1 = p_Val2_47_fu_20023_p2;

assign sext_ln856_16_fu_20178_p1 = p_Val2_50_fu_20172_p2;

assign sext_ln856_17_fu_24410_p1 = p_Val2_53_reg_41043;

assign sext_ln856_18_fu_24427_p1 = p_Val2_56_reg_41058;

assign sext_ln856_19_fu_20585_p1 = p_Val2_59_fu_20579_p2;

assign sext_ln856_1_fu_19560_p1 = p_Val2_33_reg_40614;

assign sext_ln856_20_fu_24444_p1 = p_Val2_62_reg_41073;

assign sext_ln856_21_fu_24461_p1 = p_Val2_65_reg_41088;

assign sext_ln856_22_fu_24478_p1 = p_Val2_68_reg_41103;

assign sext_ln856_23_fu_21109_p1 = p_Val2_71_reg_40965;

assign sext_ln856_24_fu_24495_p1 = p_Val2_74_reg_41118;

assign sext_ln856_25_fu_24512_p1 = p_Val2_77_reg_41133;

assign sext_ln856_26_fu_24650_p1 = p_Val2_83_reg_41191;

assign sext_ln856_27_fu_24775_p1 = p_Val2_86_reg_41222;

assign sext_ln856_28_fu_24900_p1 = p_Val2_89_reg_41253;

assign sext_ln856_29_fu_25025_p1 = p_Val2_92_reg_41284;

assign sext_ln856_2_fu_19875_p1 = p_Val2_41_reg_40687;

assign sext_ln856_30_fu_25150_p1 = p_Val2_95_reg_41315;

assign sext_ln856_31_fu_25275_p1 = p_Val2_98_reg_41346;

assign sext_ln856_32_fu_25400_p1 = p_Val2_101_reg_41377;

assign sext_ln856_33_fu_25658_p1 = p_Val2_107_fu_25652_p2;

assign sext_ln856_34_fu_25807_p1 = p_Val2_110_fu_25801_p2;

assign sext_ln856_35_fu_25956_p1 = p_Val2_113_fu_25950_p2;

assign sext_ln856_36_fu_26093_p1 = p_Val2_116_reg_41514;

assign sext_ln856_37_fu_26122_p1 = p_Val2_119_fu_26116_p2;

assign sext_ln856_38_fu_26271_p1 = p_Val2_122_fu_26265_p2;

assign sext_ln856_39_fu_26420_p1 = p_Val2_125_fu_26414_p2;

assign sext_ln856_3_fu_18489_p1 = p_Val2_2_reg_40335;

assign sext_ln856_40_fu_26569_p1 = p_Val2_128_fu_26563_p2;

assign sext_ln856_41_fu_26718_p1 = p_Val2_131_fu_26712_p2;

assign sext_ln856_42_fu_30613_p1 = p_Val2_134_reg_41756;

assign sext_ln856_43_fu_30630_p1 = p_Val2_137_reg_41783;

assign sext_ln856_44_fu_30755_p1 = p_Val2_140_reg_41814;

assign sext_ln856_45_fu_30880_p1 = p_Val2_143_reg_41845;

assign sext_ln856_46_fu_31005_p1 = p_Val2_146_reg_41876;

assign sext_ln856_47_fu_31130_p1 = p_Val2_149_reg_41907;

assign sext_ln856_48_fu_31255_p1 = p_Val2_152_reg_41926;

assign sext_ln856_49_fu_31272_p1 = p_Val2_155_reg_41953;

assign sext_ln856_4_fu_18614_p1 = p_Val2_5_reg_40366;

assign sext_ln856_50_fu_31397_p1 = p_Val2_158_reg_41972;

assign sext_ln856_51_fu_31426_p1 = p_Val2_161_fu_31420_p2;

assign sext_ln856_52_fu_31575_p1 = p_Val2_164_fu_31569_p2;

assign sext_ln856_53_fu_31724_p1 = p_Val2_167_fu_31718_p2;

assign sext_ln856_54_fu_31873_p1 = p_Val2_170_fu_31867_p2;

assign sext_ln856_55_fu_32022_p1 = p_Val2_173_fu_32016_p2;

assign sext_ln856_56_fu_32171_p1 = p_Val2_176_fu_32165_p2;

assign sext_ln856_57_fu_32320_p1 = p_Val2_179_fu_32314_p2;

assign sext_ln856_58_fu_32457_p1 = p_Val2_182_reg_42190;

assign sext_ln856_59_fu_32486_p1 = p_Val2_185_fu_32480_p2;

assign sext_ln856_5_fu_18739_p1 = p_Val2_8_reg_40385;

assign sext_ln856_60_fu_36160_p1 = p_Val2_188_reg_42398;

assign sext_ln856_61_fu_36285_p1 = p_Val2_191_reg_42429;

assign sext_ln856_62_fu_36410_p1 = p_Val2_194_reg_42460;

assign sext_ln856_63_fu_36535_p1 = p_Val2_197_reg_42491;

assign sext_ln856_64_fu_36660_p1 = p_Val2_200_reg_42522;

assign sext_ln856_65_fu_36785_p1 = p_Val2_203_reg_42541;

assign sext_ln856_66_fu_36802_p1 = p_Val2_206_reg_42568;

assign sext_ln856_67_fu_36927_p1 = p_Val2_209_reg_42599;

assign sext_ln856_68_fu_37052_p1 = p_Val2_212_reg_42630;

assign sext_ln856_69_fu_37189_p1 = p_Val2_215_fu_37183_p2;

assign sext_ln856_6_fu_18756_p1 = p_Val2_11_reg_40412;

assign sext_ln856_70_fu_37338_p1 = p_Val2_218_fu_37332_p2;

assign sext_ln856_71_fu_37487_p1 = p_Val2_221_fu_37481_p2;

assign sext_ln856_72_fu_37636_p1 = p_Val2_224_fu_37630_p2;

assign sext_ln856_73_fu_37773_p1 = p_Val2_227_reg_42765;

assign sext_ln856_74_fu_37802_p1 = p_Val2_230_fu_37796_p2;

assign sext_ln856_75_fu_37951_p1 = p_Val2_233_fu_37945_p2;

assign sext_ln856_76_fu_38100_p1 = p_Val2_236_fu_38094_p2;

assign sext_ln856_77_fu_38249_p1 = p_Val2_239_fu_38243_p2;

assign sext_ln856_7_fu_18881_p1 = p_Val2_14_reg_40443;

assign sext_ln856_8_fu_19006_p1 = p_Val2_17_reg_40474;

assign sext_ln856_9_fu_19131_p1 = p_Val2_20_reg_40493;

assign sext_ln856_fu_19543_p1 = p_Val2_31_reg_40599;

assign shl_ln1273_10_fu_33546_p3 = {{p_read_18_reg_40258_pp0_iter2_reg}, {7'd0}};

assign shl_ln1273_11_fu_33557_p3 = {{p_read_18_reg_40258_pp0_iter2_reg}, {4'd0}};

assign shl_ln1273_1_fu_18169_p1 = p_read2_int_reg;

assign shl_ln1273_1_fu_18169_p3 = {{shl_ln1273_1_fu_18169_p1}, {6'd0}};

assign shl_ln1273_2_fu_18181_p1 = p_read2_int_reg;

assign shl_ln1273_2_fu_18181_p3 = {{shl_ln1273_2_fu_18181_p1}, {2'd0}};

assign shl_ln1273_3_fu_22131_p3 = {{p_read_22_reg_40302}, {5'd0}};

assign shl_ln1273_4_fu_26876_p3 = {{p_read_21_reg_40289_pp0_iter1_reg}, {5'd0}};

assign shl_ln1273_5_fu_27384_p3 = {{p_read_21_reg_40289_pp0_iter1_reg}, {9'd0}};

assign shl_ln1273_6_fu_27401_p3 = {{p_read_21_reg_40289_pp0_iter1_reg}, {2'd0}};

assign shl_ln1273_7_fu_27662_p3 = {{p_read_21_reg_40289_pp0_iter1_reg}, {1'd0}};

assign shl_ln1273_8_fu_28173_p3 = {{p_read_20_reg_40279_pp0_iter1_reg}, {9'd0}};

assign shl_ln1273_9_fu_28184_p3 = {{p_read_20_reg_40279_pp0_iter1_reg}, {3'd0}};

assign shl_ln1273_s_fu_32960_p3 = {{p_read_19_reg_40271_pp0_iter2_reg}, {6'd0}};

assign shl_ln_fu_16411_p1 = p_read_int_reg;

assign shl_ln_fu_16411_p3 = {{shl_ln_fu_16411_p1}, {6'd0}};

assign sub_ln1273_fu_27395_p2 = ($signed(42'd0) - $signed(sext_ln1273_5_fu_27391_p1));

assign sub_ln823_1_fu_18475_p2 = (trunc_ln33_fu_16244_p1 - trunc_ln1273_1_fu_18467_p3);

assign sub_ln823_fu_16463_p2 = (trunc_ln33_1_fu_16248_p1 - trunc_ln1_fu_16427_p3);

assign tmp_105_fu_20362_p3 = r_V_15_reg_7491[32'd42];

assign tmp_111_fu_20491_p3 = r_V_16_reg_7495[32'd43];

assign tmp_117_fu_20624_p3 = r_V_17_reg_7499[32'd41];

assign tmp_123_fu_20769_p3 = r_V_18_reg_7503[32'd42];

assign tmp_129_fu_20898_p3 = r_V_19_reg_7507[32'd42];

assign tmp_12_fu_16477_p3 = sub_ln823_fu_16463_p2[32'd23];

assign tmp_135_fu_21027_p3 = r_V_20_reg_7511[32'd37];

assign tmp_138_fu_18229_p3 = r_V_21_fu_18193_p2[32'd23];

assign tmp_141_fu_18293_p3 = r_V_21_fu_18193_p2[32'd38];

assign tmp_147_fu_21173_p3 = r_V_22_reg_7515[32'd44];

assign tmp_153_fu_21302_p3 = r_V_23_reg_7519[32'd42];

assign tmp_156_fu_21434_p3 = r_V_24_fu_508_p2[32'd23];

assign tmp_159_fu_24554_p3 = r_V_24_reg_11671[32'd55];

assign tmp_15_fu_16541_p3 = r_V_2_fu_16435_p2[32'd38];

assign tmp_162_fu_21498_p3 = r_V_25_fu_497_p2[32'd23];

assign tmp_165_fu_24678_p3 = r_V_25_reg_11675[32'd43];

assign tmp_168_fu_21562_p3 = r_V_26_fu_490_p2[32'd23];

assign tmp_171_fu_24803_p3 = r_V_26_reg_11679[32'd42];

assign tmp_174_fu_21626_p3 = r_V_27_fu_541_p2[32'd23];

assign tmp_177_fu_24928_p3 = r_V_27_reg_11683[32'd43];

assign tmp_180_fu_21690_p3 = r_V_28_fu_521_p2[32'd23];

assign tmp_183_fu_25053_p3 = r_V_28_reg_11687[32'd42];

assign tmp_186_fu_21754_p3 = r_V_29_fu_538_p2[32'd23];

assign tmp_189_fu_25178_p3 = r_V_29_reg_11691[32'd40];

assign tmp_18_fu_16657_p3 = r_V_3_fu_510_p2[32'd23];

assign tmp_192_fu_21818_p3 = r_V_30_fu_488_p2[32'd23];

assign tmp_195_fu_25303_p3 = r_V_30_reg_11695[32'd40];

assign tmp_198_fu_21882_p3 = r_V_31_fu_496_p2[32'd23];

assign tmp_201_fu_25428_p3 = r_V_31_reg_11699[32'd45];

assign tmp_204_fu_21942_p3 = r_V_32_fu_499_p2[32'd23];

assign tmp_207_fu_25550_p3 = r_V_32_reg_11703[32'd55];

assign tmp_213_fu_25697_p3 = r_V_33_reg_11707[32'd50];

assign tmp_219_fu_25846_p3 = r_V_34_reg_11711[32'd43];

assign tmp_21_fu_18784_p3 = r_V_3_reg_7447[32'd44];

assign tmp_225_fu_25995_p3 = r_V_35_reg_11715[32'd41];

assign tmp_228_fu_22178_p3 = r_V_36_fu_22142_p2[32'd23];

assign tmp_231_fu_22242_p3 = r_V_36_fu_22142_p2[32'd37];

assign tmp_237_fu_26161_p3 = r_V_37_reg_11719[32'd42];

assign tmp_243_fu_26310_p3 = r_V_38_reg_11723[32'd43];

assign tmp_249_fu_26459_p3 = r_V_39_reg_11727[32'd42];

assign tmp_24_fu_16721_p3 = r_V_4_fu_526_p2[32'd23];

assign tmp_255_fu_26608_p3 = r_V_40_reg_11731[32'd44];

assign tmp_261_fu_26757_p3 = r_V_41_reg_11735[32'd52];

assign tmp_267_fu_26978_p3 = r_V_42_fu_26887_p2[32'd37];

assign tmp_270_fu_27094_p3 = r_V_43_fu_531_p2[32'd23];

assign tmp_273_fu_30658_p3 = r_V_43_reg_14203[32'd42];

assign tmp_276_fu_27158_p3 = r_V_44_fu_520_p2[32'd23];

assign tmp_279_fu_30783_p3 = r_V_44_reg_14207[32'd41];

assign tmp_27_fu_18909_p3 = r_V_4_reg_7451[32'd42];

assign tmp_282_fu_27222_p3 = r_V_45_fu_506_p2[32'd23];

assign tmp_285_fu_30908_p3 = r_V_45_reg_14211[32'd44];

assign tmp_288_fu_27286_p3 = r_V_46_fu_530_p2[32'd23];

assign tmp_291_fu_31033_p3 = r_V_46_reg_14215[32'd43];

assign tmp_294_fu_27350_p3 = r_V_47_fu_471_p2[32'd23];

assign tmp_297_fu_31158_p3 = r_V_47_reg_14219[32'd42];

assign tmp_300_fu_27448_p3 = r_V_48_fu_27412_p2[32'd23];

assign tmp_303_fu_27512_p3 = r_V_48_fu_27412_p2[32'd41];

assign tmp_306_fu_27628_p3 = r_V_49_fu_480_p2[32'd23];

assign tmp_309_fu_31300_p3 = r_V_49_reg_14223[32'd42];

assign tmp_30_fu_16785_p3 = r_V_5_fu_500_p2[32'd23];

assign tmp_312_fu_27709_p3 = r_V_50_fu_27673_p2[32'd23];

assign tmp_315_fu_27773_p3 = r_V_50_fu_27673_p2[32'd41];

assign tmp_321_fu_31465_p3 = r_V_51_reg_14227[32'd42];

assign tmp_327_fu_31614_p3 = r_V_52_reg_14231[32'd41];

assign tmp_333_fu_31763_p3 = r_V_53_reg_14235[32'd43];

assign tmp_339_fu_31912_p3 = r_V_54_reg_14239[32'd44];

assign tmp_33_fu_19034_p3 = r_V_5_reg_7455[32'd42];

assign tmp_345_fu_32061_p3 = r_V_55_reg_14243[32'd44];

assign tmp_351_fu_32210_p3 = r_V_56_reg_14247[32'd43];

assign tmp_357_fu_32359_p3 = r_V_57_reg_14251[32'd44];

assign tmp_360_fu_28231_p3 = r_V_58_fu_28195_p2[32'd23];

assign tmp_363_fu_28295_p3 = r_V_58_fu_28195_p2[32'd41];

assign tmp_369_fu_32525_p3 = r_V_59_reg_14255[32'd43];

assign tmp_36_fu_16855_p3 = r_V_6_fu_16819_p2[32'd23];

assign tmp_372_fu_32670_p3 = r_V_60_fu_474_p2[32'd23];

assign tmp_375_fu_36188_p3 = r_V_60_reg_16179[32'd41];

assign tmp_378_fu_32734_p3 = r_V_61_fu_543_p2[32'd23];

assign tmp_381_fu_36313_p3 = r_V_61_reg_16183[32'd42];

assign tmp_384_fu_32798_p3 = r_V_62_fu_477_p2[32'd23];

assign tmp_387_fu_36438_p3 = r_V_62_reg_16187[32'd43];

assign tmp_390_fu_32862_p3 = r_V_63_fu_545_p2[32'd23];

assign tmp_393_fu_36563_p3 = r_V_63_reg_16191[32'd41];

assign tmp_396_fu_32926_p3 = r_V_64_fu_533_p2[32'd23];

assign tmp_399_fu_36688_p3 = r_V_64_reg_16195[32'd43];

assign tmp_39_fu_16919_p3 = r_V_6_fu_16819_p2[32'd38];

assign tmp_3_fu_18517_p3 = r_V_reg_7439[32'd46];

assign tmp_402_fu_33007_p3 = r_V_65_fu_32971_p2[32'd23];

assign tmp_405_fu_33071_p3 = r_V_65_fu_32971_p2[32'd38];

assign tmp_408_fu_33187_p3 = r_V_66_fu_511_p2[32'd23];

assign tmp_411_fu_36830_p3 = r_V_66_reg_16199[32'd42];

assign tmp_414_fu_33251_p3 = r_V_67_fu_522_p2[32'd23];

assign tmp_417_fu_36955_p3 = r_V_67_reg_16203[32'd43];

assign tmp_420_fu_33315_p3 = r_V_68_fu_544_p2[32'd23];

assign tmp_423_fu_37080_p3 = r_V_68_reg_16207[32'd41];

assign tmp_429_fu_37228_p3 = r_V_69_reg_16211[32'd43];

assign tmp_42_fu_17031_p3 = r_V_7_fu_537_p2[32'd23];

assign tmp_435_fu_37377_p3 = r_V_70_reg_16215[32'd42];

assign tmp_441_fu_37526_p3 = r_V_71_reg_16219[32'd41];

assign tmp_447_fu_37675_p3 = r_V_72_reg_16223[32'd42];

assign tmp_450_fu_33604_p3 = r_V_73_fu_33568_p2[32'd23];

assign tmp_453_fu_33668_p3 = r_V_73_fu_33568_p2[32'd39];

assign tmp_459_fu_37841_p3 = r_V_74_reg_16227[32'd40];

assign tmp_45_fu_19173_p3 = r_V_7_reg_7459[32'd56];

assign tmp_465_fu_37990_p3 = r_V_75_reg_16231[32'd39];

assign tmp_471_fu_38139_p3 = r_V_76_reg_16235[32'd45];

assign tmp_477_fu_38288_p3 = r_V_77_reg_16239[32'd53];

assign tmp_48_fu_17095_p3 = r_V_8_fu_514_p2[32'd23];

assign tmp_51_fu_19297_p3 = r_V_8_reg_7463[32'd44];

assign tmp_57_fu_19445_p3 = r_V_9_reg_7467[32'd42];

assign tmp_60_fu_17219_p1 = p_read1_int_reg;

assign tmp_60_fu_17219_p3 = tmp_60_fu_17219_p1[32'd14];

assign tmp_63_fu_17271_p1 = p_read1_int_reg;

assign tmp_63_fu_17271_p3 = tmp_63_fu_17271_p1[32'd31];

assign tmp_65_fu_17391_p1 = p_read1_int_reg;

assign tmp_65_fu_17391_p3 = tmp_65_fu_17391_p1[32'd18];

assign tmp_6_fu_16377_p3 = r_V_1_fu_470_p2[32'd23];

assign tmp_72_fu_19628_p3 = r_V_10_reg_7471[32'd44];

assign tmp_78_fu_19777_p3 = r_V_11_reg_7475[32'd44];

assign tmp_80_fu_17619_p1 = p_read1_int_reg;

assign tmp_80_fu_17619_p3 = tmp_80_fu_17619_p1[32'd15];

assign tmp_84_fu_17771_p3 = r_V_12_fu_489_p2[32'd23];

assign tmp_87_fu_19920_p3 = r_V_12_reg_7479[32'd41];

assign tmp_93_fu_20068_p3 = r_V_13_reg_7483[32'd42];

assign tmp_99_fu_20217_p3 = r_V_14_reg_7487[32'd44];

assign tmp_9_fu_18642_p3 = r_V_1_reg_7443[32'd41];

assign tmp_fu_16313_p3 = r_V_fu_519_p2[32'd23];

assign trunc_ln1273_1_fu_18467_p3 = {{trunc_ln1273_2_fu_18463_p1}, {5'd0}};

assign trunc_ln1273_2_fu_18463_p0 = p_read5_int_reg;

assign trunc_ln1273_2_fu_18463_p1 = trunc_ln1273_2_fu_18463_p0[18:0];

assign trunc_ln1273_fu_16423_p0 = p_read_int_reg;

assign trunc_ln1273_fu_16423_p1 = trunc_ln1273_fu_16423_p0[17:0];

assign trunc_ln1_fu_16427_p3 = {{trunc_ln1273_fu_16423_p1}, {6'd0}};

assign trunc_ln33_1_fu_16248_p0 = p_read_int_reg;

assign trunc_ln33_1_fu_16248_p1 = trunc_ln33_1_fu_16248_p0[23:0];

assign trunc_ln33_fu_16244_p0 = p_read5_int_reg;

assign trunc_ln33_fu_16244_p1 = trunc_ln33_fu_16244_p0[23:0];

assign underflow_100_fu_28575_p2 = (xor_ln896_181_fu_28569_p2 & p_Result_279_fu_28536_p3);

assign underflow_101_fu_28638_p2 = (xor_ln896_182_fu_28633_p2 & p_Result_281_reg_41716);

assign underflow_102_fu_28733_p2 = (xor_ln896_183_fu_28727_p2 & p_Result_283_fu_28694_p3);

assign underflow_103_fu_28833_p2 = (xor_ln896_184_fu_28827_p2 & p_Result_285_fu_28794_p3);

assign underflow_104_fu_28933_p2 = (xor_ln896_185_fu_28927_p2 & p_Result_287_fu_28894_p3);

assign underflow_105_fu_28996_p2 = (xor_ln896_186_fu_28991_p2 & p_Result_289_reg_41736);

assign underflow_106_fu_29091_p2 = (xor_ln896_187_fu_29085_p2 & p_Result_291_fu_29052_p3);

assign underflow_107_fu_29191_p2 = (xor_ln896_188_fu_29185_p2 & p_Result_293_fu_29152_p3);

assign underflow_108_fu_29293_p2 = (xor_ln896_189_fu_29287_p2 & p_Result_295_fu_29253_p3);

assign underflow_109_fu_29395_p2 = (xor_ln896_190_fu_29389_p2 & p_Result_297_fu_29355_p3);

assign underflow_10_fu_17357_p2 = (xor_ln896_253_fu_17351_p2 & p_Result_30_fu_17189_p3);

assign underflow_110_fu_29497_p2 = (xor_ln896_191_fu_29491_p2 & p_Result_299_fu_29457_p3);

assign underflow_111_fu_29599_p2 = (xor_ln896_192_fu_29593_p2 & p_Result_301_fu_29559_p3);

assign underflow_112_fu_29701_p2 = (xor_ln896_193_fu_29695_p2 & p_Result_303_fu_29661_p3);

assign underflow_113_fu_29803_p2 = (xor_ln896_194_fu_29797_p2 & p_Result_305_fu_29763_p3);

assign underflow_114_fu_29905_p2 = (xor_ln896_195_fu_29899_p2 & p_Result_307_fu_29865_p3);

assign underflow_115_fu_30007_p2 = (xor_ln896_196_fu_30001_p2 & p_Result_309_fu_29967_p3);

assign underflow_116_fu_30109_p2 = (xor_ln896_197_fu_30103_p2 & p_Result_311_fu_30069_p3);

assign underflow_117_fu_33937_p2 = (xor_ln896_198_fu_33932_p2 & p_Result_313_reg_42234);

assign underflow_118_fu_33995_p2 = (xor_ln896_199_fu_33990_p2 & p_Result_315_reg_42254);

assign underflow_119_fu_30283_p2 = (xor_ln896_200_fu_30277_p2 & p_Result_317_fu_30243_p3);

assign underflow_11_fu_17501_p2 = (xor_ln896_254_fu_17495_p2 & p_Result_30_fu_17189_p3);

assign underflow_120_fu_34053_p2 = (xor_ln896_201_fu_34048_p2 & p_Result_319_reg_42280);

assign underflow_121_fu_34111_p2 = (xor_ln896_202_fu_34106_p2 & p_Result_321_reg_42300);

assign underflow_122_fu_34169_p2 = (xor_ln896_203_fu_34164_p2 & p_Result_323_reg_42320);

assign underflow_123_fu_30493_p2 = (xor_ln896_204_fu_30487_p2 & p_Result_325_fu_30453_p3);

assign underflow_124_fu_34227_p2 = (xor_ln896_205_fu_34222_p2 & p_Result_327_reg_42346);

assign underflow_125_fu_34285_p2 = (xor_ln896_206_fu_34280_p2 & p_Result_329_reg_42366);

assign underflow_126_fu_34382_p2 = (xor_ln896_207_fu_34376_p2 & p_Result_331_fu_34342_p3);

assign underflow_127_fu_34484_p2 = (xor_ln896_208_fu_34478_p2 & p_Result_333_fu_34444_p3);

assign underflow_128_fu_34584_p2 = (xor_ln896_209_fu_34578_p2 & p_Result_335_fu_34545_p3);

assign underflow_129_fu_34686_p2 = (xor_ln896_210_fu_34680_p2 & p_Result_337_fu_34646_p3);

assign underflow_12_fu_19699_p2 = (xor_ln896_255_fu_19693_p2 & p_Result_35_reg_40629);

assign underflow_130_fu_34788_p2 = (xor_ln896_211_fu_34782_p2 & p_Result_339_fu_34748_p3);

assign underflow_131_fu_34890_p2 = (xor_ln896_212_fu_34884_p2 & p_Result_341_fu_34850_p3);

assign underflow_132_fu_34990_p2 = (xor_ln896_213_fu_34984_p2 & p_Result_343_fu_34951_p3);

assign underflow_133_fu_35092_p2 = (xor_ln896_214_fu_35086_p2 & p_Result_345_fu_35052_p3);

assign underflow_134_fu_35194_p2 = (xor_ln896_215_fu_35188_p2 & p_Result_347_fu_35154_p3);

assign underflow_135_fu_35296_p2 = (xor_ln896_216_fu_35290_p2 & p_Result_349_fu_35256_p3);

assign underflow_136_fu_35398_p2 = (xor_ln896_217_fu_35392_p2 & p_Result_351_fu_35358_p3);

assign underflow_137_fu_35500_p2 = (xor_ln896_218_fu_35494_p2 & p_Result_353_fu_35460_p3);

assign underflow_138_fu_35602_p2 = (xor_ln896_219_fu_35596_p2 & p_Result_355_fu_35562_p3);

assign underflow_139_fu_35704_p2 = (xor_ln896_220_fu_35698_p2 & p_Result_357_fu_35664_p3);

assign underflow_13_fu_19848_p2 = (xor_ln896_256_fu_19842_p2 & p_Result_38_reg_40658);

assign underflow_140_fu_35806_p2 = (xor_ln896_221_fu_35800_p2 & p_Result_359_fu_35766_p3);

assign underflow_141_fu_35908_p2 = (xor_ln896_222_fu_35902_p2 & p_Result_361_fu_35868_p3);

assign underflow_142_fu_36010_p2 = (xor_ln896_223_fu_36004_p2 & p_Result_363_fu_35970_p3);

assign underflow_143_fu_36112_p2 = (xor_ln896_224_fu_36106_p2 & p_Result_365_fu_36072_p3);

assign underflow_144_fu_38438_p2 = (xor_ln896_225_fu_38432_p2 & p_Result_367_fu_38399_p3);

assign underflow_145_fu_38538_p2 = (xor_ln896_226_fu_38532_p2 & p_Result_369_fu_38499_p3);

assign underflow_146_fu_38638_p2 = (xor_ln896_227_fu_38632_p2 & p_Result_371_fu_38599_p3);

assign underflow_147_fu_38738_p2 = (xor_ln896_228_fu_38732_p2 & p_Result_373_fu_38699_p3);

assign underflow_148_fu_38838_p2 = (xor_ln896_229_fu_38832_p2 & p_Result_375_fu_38799_p3);

assign underflow_149_fu_38938_p2 = (xor_ln896_230_fu_38932_p2 & p_Result_377_fu_38899_p3);

assign underflow_14_fu_17729_p2 = (xor_ln896_257_fu_17723_p2 & p_Result_30_fu_17189_p3);

assign underflow_150_fu_39038_p2 = (xor_ln896_231_fu_39032_p2 & p_Result_379_fu_38999_p3);

assign underflow_151_fu_39138_p2 = (xor_ln896_232_fu_39132_p2 & p_Result_381_fu_39099_p3);

assign underflow_152_fu_39238_p2 = (xor_ln896_233_fu_39232_p2 & p_Result_383_fu_39199_p3);

assign underflow_153_fu_39340_p2 = (xor_ln896_234_fu_39334_p2 & p_Result_385_fu_39300_p3);

assign underflow_154_fu_39442_p2 = (xor_ln896_235_fu_39436_p2 & p_Result_387_fu_39402_p3);

assign underflow_155_fu_39544_p2 = (xor_ln896_236_fu_39538_p2 & p_Result_389_fu_39504_p3);

assign underflow_156_fu_39646_p2 = (xor_ln896_237_fu_39640_p2 & p_Result_391_fu_39606_p3);

assign underflow_157_fu_39748_p2 = (xor_ln896_238_fu_39742_p2 & p_Result_393_fu_39708_p3);

assign underflow_158_fu_39850_p2 = (xor_ln896_239_fu_39844_p2 & p_Result_395_fu_39810_p3);

assign underflow_159_fu_39952_p2 = (xor_ln896_240_fu_39946_p2 & p_Result_397_fu_39912_p3);

assign underflow_15_fu_19990_p2 = (xor_ln896_258_fu_19984_p2 & p_Result_43_reg_40702);

assign underflow_160_fu_40054_p2 = (xor_ln896_241_fu_40048_p2 & p_Result_399_fu_40014_p3);

assign underflow_161_fu_40156_p2 = (xor_ln896_242_fu_40150_p2 & p_Result_401_fu_40116_p3);

assign underflow_16_fu_20139_p2 = (xor_ln896_259_fu_20133_p2 & p_Result_46_reg_40733);

assign underflow_17_fu_20288_p2 = (xor_ln896_260_fu_20282_p2 & p_Result_49_reg_40762);

assign underflow_18_fu_20433_p2 = (xor_ln896_261_fu_20427_p2 & p_Result_52_reg_40791);

assign underflow_19_fu_20562_p2 = (xor_ln896_262_fu_20556_p2 & p_Result_55_reg_40820);

assign underflow_1_fu_18712_p2 = (xor_ln896_244_fu_18706_p2 & p_Result_3_reg_40354);

assign underflow_20_fu_20695_p2 = (xor_ln896_263_fu_20689_p2 & p_Result_58_reg_40849);

assign underflow_21_fu_20840_p2 = (xor_ln896_264_fu_20834_p2 & p_Result_61_reg_40878);

assign underflow_22_fu_20969_p2 = (xor_ln896_265_fu_20963_p2 & p_Result_64_reg_40907);

assign underflow_23_fu_21098_p2 = (xor_ln896_266_fu_21092_p2 & p_Result_67_reg_40936);

assign underflow_24_fu_18367_p2 = (xor_ln896_267_fu_18361_p2 & p_Result_70_fu_18199_p3);

assign underflow_25_fu_21244_p2 = (xor_ln896_268_fu_21238_p2 & p_Result_73_reg_40980);

assign underflow_26_fu_21373_p2 = (xor_ln896_269_fu_21367_p2 & p_Result_76_reg_41009);

assign underflow_27_fu_24624_p2 = (xor_ln896_270_fu_24618_p2 & p_Result_79_reg_41148);

assign underflow_28_fu_24748_p2 = (xor_ln896_271_fu_24742_p2 & p_Result_82_reg_41179);

assign underflow_29_fu_24873_p2 = (xor_ln896_272_fu_24867_p2 & p_Result_85_reg_41210);

assign underflow_2_fu_16615_p2 = (xor_ln896_245_fu_16609_p2 & p_Result_6_fu_16441_p3);

assign underflow_30_fu_24998_p2 = (xor_ln896_273_fu_24992_p2 & p_Result_88_reg_41241);

assign underflow_31_fu_25123_p2 = (xor_ln896_274_fu_25117_p2 & p_Result_91_reg_41272);

assign underflow_32_fu_25248_p2 = (xor_ln896_275_fu_25242_p2 & p_Result_94_reg_41303);

assign underflow_33_fu_25373_p2 = (xor_ln896_276_fu_25367_p2 & p_Result_97_reg_41334);

assign underflow_34_fu_25498_p2 = (xor_ln896_277_fu_25492_p2 & p_Result_100_reg_41365);

assign underflow_35_fu_25620_p2 = (xor_ln896_278_fu_25614_p2 & p_Result_103_reg_41396);

assign underflow_36_fu_25768_p2 = (xor_ln896_279_fu_25762_p2 & p_Result_106_reg_41427);

assign underflow_37_fu_25917_p2 = (xor_ln896_280_fu_25911_p2 & p_Result_109_reg_41456);

assign underflow_38_fu_26066_p2 = (xor_ln896_281_fu_26060_p2 & p_Result_112_reg_41485);

assign underflow_39_fu_22316_p2 = (xor_ln896_282_fu_22310_p2 & p_Result_115_fu_22148_p3);

assign underflow_3_fu_18854_p2 = (xor_ln896_246_fu_18848_p2 & p_Result_9_reg_40400);

assign underflow_40_fu_26232_p2 = (xor_ln896_283_fu_26226_p2 & p_Result_118_reg_41529);

assign underflow_41_fu_26381_p2 = (xor_ln896_284_fu_26375_p2 & p_Result_121_reg_41558);

assign underflow_42_fu_26530_p2 = (xor_ln896_285_fu_26524_p2 & p_Result_124_reg_41587);

assign underflow_43_fu_26679_p2 = (xor_ln896_286_fu_26673_p2 & p_Result_127_reg_41616);

assign underflow_44_fu_26828_p2 = (xor_ln896_287_fu_26822_p2 & p_Result_130_reg_41645);

assign underflow_45_fu_27052_p2 = (xor_ln896_288_fu_27046_p2 & p_Result_133_fu_26893_p3);

assign underflow_46_fu_30728_p2 = (xor_ln896_289_fu_30722_p2 & p_Result_136_reg_41771);

assign underflow_47_fu_30853_p2 = (xor_ln896_290_fu_30847_p2 & p_Result_139_reg_41802);

assign underflow_48_fu_30978_p2 = (xor_ln896_291_fu_30972_p2 & p_Result_142_reg_41833);

assign underflow_49_fu_31103_p2 = (xor_ln896_292_fu_31097_p2 & p_Result_145_reg_41864);

assign underflow_4_fu_18979_p2 = (xor_ln896_247_fu_18973_p2 & p_Result_12_reg_40431);

assign underflow_50_fu_31228_p2 = (xor_ln896_293_fu_31222_p2 & p_Result_148_reg_41895);

assign underflow_51_fu_27586_p2 = (xor_ln896_294_fu_27580_p2 & p_Result_151_fu_27418_p3);

assign underflow_52_fu_31370_p2 = (xor_ln896_295_fu_31364_p2 & p_Result_154_reg_41941);

assign underflow_53_fu_27847_p2 = (xor_ln896_296_fu_27841_p2 & p_Result_157_fu_27679_p3);

assign underflow_54_fu_31536_p2 = (xor_ln896_297_fu_31530_p2 & p_Result_160_reg_41987);

assign underflow_55_fu_31685_p2 = (xor_ln896_298_fu_31679_p2 & p_Result_163_reg_42016);

assign underflow_56_fu_31834_p2 = (xor_ln896_299_fu_31828_p2 & p_Result_166_reg_42045);

assign underflow_57_fu_31983_p2 = (xor_ln896_300_fu_31977_p2 & p_Result_169_reg_42074);

assign underflow_58_fu_32132_p2 = (xor_ln896_301_fu_32126_p2 & p_Result_172_reg_42103);

assign underflow_59_fu_32281_p2 = (xor_ln896_302_fu_32275_p2 & p_Result_175_reg_42132);

assign underflow_5_fu_19104_p2 = (xor_ln896_248_fu_19098_p2 & p_Result_15_reg_40462);

assign underflow_60_fu_32430_p2 = (xor_ln896_303_fu_32424_p2 & p_Result_178_reg_42161);

assign underflow_61_fu_28369_p2 = (xor_ln896_304_fu_28363_p2 & p_Result_181_fu_28201_p3);

assign underflow_62_fu_32596_p2 = (xor_ln896_305_fu_32590_p2 & p_Result_184_reg_42205);

assign underflow_63_fu_36258_p2 = (xor_ln896_306_fu_36252_p2 & p_Result_187_reg_42386);

assign underflow_64_fu_36383_p2 = (xor_ln896_307_fu_36377_p2 & p_Result_190_reg_42417);

assign underflow_65_fu_36508_p2 = (xor_ln896_308_fu_36502_p2 & p_Result_193_reg_42448);

assign underflow_66_fu_36633_p2 = (xor_ln896_309_fu_36627_p2 & p_Result_196_reg_42479);

assign underflow_67_fu_36758_p2 = (xor_ln896_310_fu_36752_p2 & p_Result_199_reg_42510);

assign underflow_68_fu_33145_p2 = (xor_ln896_311_fu_33139_p2 & p_Result_202_fu_32977_p3);

assign underflow_69_fu_36900_p2 = (xor_ln896_312_fu_36894_p2 & p_Result_205_reg_42556);

assign underflow_6_fu_16993_p2 = (xor_ln896_249_fu_16987_p2 & p_Result_18_fu_16825_p3);

assign underflow_70_fu_37025_p2 = (xor_ln896_313_fu_37019_p2 & p_Result_208_reg_42587);

assign underflow_71_fu_37150_p2 = (xor_ln896_314_fu_37144_p2 & p_Result_211_reg_42618);

assign underflow_72_fu_37299_p2 = (xor_ln896_315_fu_37293_p2 & p_Result_214_reg_42649);

assign underflow_73_fu_37448_p2 = (xor_ln896_316_fu_37442_p2 & p_Result_217_reg_42678);

assign underflow_74_fu_37597_p2 = (xor_ln896_317_fu_37591_p2 & p_Result_220_reg_42707);

assign underflow_75_fu_37746_p2 = (xor_ln896_318_fu_37740_p2 & p_Result_223_reg_42736);

assign underflow_76_fu_33742_p2 = (xor_ln896_319_fu_33736_p2 & p_Result_226_fu_33574_p3);

assign underflow_77_fu_37912_p2 = (xor_ln896_320_fu_37906_p2 & p_Result_229_reg_42780);

assign underflow_78_fu_38061_p2 = (xor_ln896_321_fu_38055_p2 & p_Result_232_reg_42809);

assign underflow_79_fu_38210_p2 = (xor_ln896_322_fu_38204_p2 & p_Result_235_reg_42838);

assign underflow_7_fu_19243_p2 = (xor_ln896_250_fu_19237_p2 & p_Result_21_reg_40508);

assign underflow_80_fu_38359_p2 = (xor_ln896_323_fu_38353_p2 & p_Result_238_reg_42867);

assign underflow_81_fu_22588_p2 = (xor_ln896_162_fu_22582_p2 & p_Result_241_fu_22548_p3);

assign underflow_82_fu_22686_p2 = (xor_ln896_163_fu_22680_p2 & p_Result_243_fu_22646_p3);

assign underflow_83_fu_22784_p2 = (xor_ln896_164_fu_22778_p2 & p_Result_245_fu_22744_p3);

assign underflow_84_fu_22882_p2 = (xor_ln896_165_fu_22876_p2 & p_Result_247_fu_22842_p3);

assign underflow_85_fu_22980_p2 = (xor_ln896_166_fu_22974_p2 & p_Result_249_fu_22940_p3);

assign underflow_86_fu_23078_p2 = (xor_ln896_167_fu_23072_p2 & p_Result_251_fu_23038_p3);

assign underflow_87_fu_23176_p2 = (xor_ln896_168_fu_23170_p2 & p_Result_253_fu_23136_p3);

assign underflow_88_fu_23274_p2 = (xor_ln896_169_fu_23268_p2 & p_Result_255_fu_23234_p3);

assign underflow_89_fu_23372_p2 = (xor_ln896_170_fu_23366_p2 & p_Result_257_fu_23332_p3);

assign underflow_8_fu_19367_p2 = (xor_ln896_251_fu_19361_p2 & p_Result_24_reg_40539);

assign underflow_90_fu_23474_p2 = (xor_ln896_171_fu_23468_p2 & p_Result_259_fu_23434_p3);

assign underflow_91_fu_23576_p2 = (xor_ln896_172_fu_23570_p2 & p_Result_261_fu_23536_p3);

assign underflow_92_fu_23678_p2 = (xor_ln896_173_fu_23672_p2 & p_Result_263_fu_23638_p3);

assign underflow_93_fu_23780_p2 = (xor_ln896_174_fu_23774_p2 & p_Result_265_fu_23740_p3);

assign underflow_94_fu_23882_p2 = (xor_ln896_175_fu_23876_p2 & p_Result_267_fu_23842_p3);

assign underflow_95_fu_23984_p2 = (xor_ln896_176_fu_23978_p2 & p_Result_269_fu_23944_p3);

assign underflow_96_fu_24086_p2 = (xor_ln896_177_fu_24080_p2 & p_Result_271_fu_24046_p3);

assign underflow_97_fu_24188_p2 = (xor_ln896_178_fu_24182_p2 & p_Result_273_fu_24148_p3);

assign underflow_98_fu_24290_p2 = (xor_ln896_179_fu_24284_p2 & p_Result_275_fu_24250_p3);

assign underflow_99_fu_28475_p2 = (xor_ln896_180_fu_28469_p2 & p_Result_277_fu_28436_p3);

assign underflow_9_fu_19516_p2 = (xor_ln896_252_fu_19510_p2 & p_Result_27_reg_40570);

assign underflow_fu_18587_p2 = (xor_ln896_243_fu_18581_p2 & p_Result_s_reg_40323);

assign xor_ln302_100_fu_34896_p2 = (p_Result_342_fu_34864_p3 ^ p_Result_341_fu_34850_p3);

assign xor_ln302_101_fu_34902_p2 = (xor_ln302_100_fu_34896_p2 ^ 1'd1);

assign xor_ln302_102_fu_34996_p2 = (p_Result_344_fu_34964_p3 ^ p_Result_343_fu_34951_p3);

assign xor_ln302_103_fu_35002_p2 = (xor_ln302_102_fu_34996_p2 ^ 1'd1);

assign xor_ln302_104_fu_35098_p2 = (p_Result_346_fu_35066_p3 ^ p_Result_345_fu_35052_p3);

assign xor_ln302_105_fu_35104_p2 = (xor_ln302_104_fu_35098_p2 ^ 1'd1);

assign xor_ln302_106_fu_35200_p2 = (p_Result_348_fu_35168_p3 ^ p_Result_347_fu_35154_p3);

assign xor_ln302_107_fu_35206_p2 = (xor_ln302_106_fu_35200_p2 ^ 1'd1);

assign xor_ln302_108_fu_35302_p2 = (p_Result_350_fu_35270_p3 ^ p_Result_349_fu_35256_p3);

assign xor_ln302_109_fu_35308_p2 = (xor_ln302_108_fu_35302_p2 ^ 1'd1);

assign xor_ln302_10_fu_23084_p2 = (p_Result_252_fu_23052_p3 ^ p_Result_251_fu_23038_p3);

assign xor_ln302_110_fu_35404_p2 = (p_Result_352_fu_35372_p3 ^ p_Result_351_fu_35358_p3);

assign xor_ln302_111_fu_35410_p2 = (xor_ln302_110_fu_35404_p2 ^ 1'd1);

assign xor_ln302_112_fu_35506_p2 = (p_Result_354_fu_35474_p3 ^ p_Result_353_fu_35460_p3);

assign xor_ln302_113_fu_35512_p2 = (xor_ln302_112_fu_35506_p2 ^ 1'd1);

assign xor_ln302_114_fu_35608_p2 = (p_Result_356_fu_35576_p3 ^ p_Result_355_fu_35562_p3);

assign xor_ln302_115_fu_35614_p2 = (xor_ln302_114_fu_35608_p2 ^ 1'd1);

assign xor_ln302_116_fu_35710_p2 = (p_Result_358_fu_35678_p3 ^ p_Result_357_fu_35664_p3);

assign xor_ln302_117_fu_35716_p2 = (xor_ln302_116_fu_35710_p2 ^ 1'd1);

assign xor_ln302_118_fu_35812_p2 = (p_Result_360_fu_35780_p3 ^ p_Result_359_fu_35766_p3);

assign xor_ln302_119_fu_35818_p2 = (xor_ln302_118_fu_35812_p2 ^ 1'd1);

assign xor_ln302_11_fu_23090_p2 = (xor_ln302_10_fu_23084_p2 ^ 1'd1);

assign xor_ln302_120_fu_35914_p2 = (p_Result_362_fu_35882_p3 ^ p_Result_361_fu_35868_p3);

assign xor_ln302_121_fu_35920_p2 = (xor_ln302_120_fu_35914_p2 ^ 1'd1);

assign xor_ln302_122_fu_36016_p2 = (p_Result_364_fu_35984_p3 ^ p_Result_363_fu_35970_p3);

assign xor_ln302_123_fu_36022_p2 = (xor_ln302_122_fu_36016_p2 ^ 1'd1);

assign xor_ln302_124_fu_36118_p2 = (p_Result_366_fu_36086_p3 ^ p_Result_365_fu_36072_p3);

assign xor_ln302_125_fu_36124_p2 = (xor_ln302_124_fu_36118_p2 ^ 1'd1);

assign xor_ln302_126_fu_38444_p2 = (p_Result_368_fu_38412_p3 ^ p_Result_367_fu_38399_p3);

assign xor_ln302_127_fu_38450_p2 = (xor_ln302_126_fu_38444_p2 ^ 1'd1);

assign xor_ln302_128_fu_38544_p2 = (p_Result_370_fu_38512_p3 ^ p_Result_369_fu_38499_p3);

assign xor_ln302_129_fu_38550_p2 = (xor_ln302_128_fu_38544_p2 ^ 1'd1);

assign xor_ln302_12_fu_23182_p2 = (p_Result_254_fu_23150_p3 ^ p_Result_253_fu_23136_p3);

assign xor_ln302_130_fu_38644_p2 = (p_Result_372_fu_38612_p3 ^ p_Result_371_fu_38599_p3);

assign xor_ln302_131_fu_38650_p2 = (xor_ln302_130_fu_38644_p2 ^ 1'd1);

assign xor_ln302_132_fu_38744_p2 = (p_Result_374_fu_38712_p3 ^ p_Result_373_fu_38699_p3);

assign xor_ln302_133_fu_38750_p2 = (xor_ln302_132_fu_38744_p2 ^ 1'd1);

assign xor_ln302_134_fu_38844_p2 = (p_Result_376_fu_38812_p3 ^ p_Result_375_fu_38799_p3);

assign xor_ln302_135_fu_38850_p2 = (xor_ln302_134_fu_38844_p2 ^ 1'd1);

assign xor_ln302_136_fu_38944_p2 = (p_Result_378_fu_38912_p3 ^ p_Result_377_fu_38899_p3);

assign xor_ln302_137_fu_38950_p2 = (xor_ln302_136_fu_38944_p2 ^ 1'd1);

assign xor_ln302_138_fu_39044_p2 = (p_Result_380_fu_39012_p3 ^ p_Result_379_fu_38999_p3);

assign xor_ln302_139_fu_39050_p2 = (xor_ln302_138_fu_39044_p2 ^ 1'd1);

assign xor_ln302_13_fu_23188_p2 = (xor_ln302_12_fu_23182_p2 ^ 1'd1);

assign xor_ln302_140_fu_39144_p2 = (p_Result_382_fu_39112_p3 ^ p_Result_381_fu_39099_p3);

assign xor_ln302_141_fu_39150_p2 = (xor_ln302_140_fu_39144_p2 ^ 1'd1);

assign xor_ln302_142_fu_39244_p2 = (p_Result_384_fu_39212_p3 ^ p_Result_383_fu_39199_p3);

assign xor_ln302_143_fu_39250_p2 = (xor_ln302_142_fu_39244_p2 ^ 1'd1);

assign xor_ln302_144_fu_39346_p2 = (p_Result_386_fu_39314_p3 ^ p_Result_385_fu_39300_p3);

assign xor_ln302_145_fu_39352_p2 = (xor_ln302_144_fu_39346_p2 ^ 1'd1);

assign xor_ln302_146_fu_39448_p2 = (p_Result_388_fu_39416_p3 ^ p_Result_387_fu_39402_p3);

assign xor_ln302_147_fu_39454_p2 = (xor_ln302_146_fu_39448_p2 ^ 1'd1);

assign xor_ln302_148_fu_39550_p2 = (p_Result_390_fu_39518_p3 ^ p_Result_389_fu_39504_p3);

assign xor_ln302_149_fu_39556_p2 = (xor_ln302_148_fu_39550_p2 ^ 1'd1);

assign xor_ln302_14_fu_23280_p2 = (p_Result_256_fu_23248_p3 ^ p_Result_255_fu_23234_p3);

assign xor_ln302_150_fu_39652_p2 = (p_Result_392_fu_39620_p3 ^ p_Result_391_fu_39606_p3);

assign xor_ln302_151_fu_39658_p2 = (xor_ln302_150_fu_39652_p2 ^ 1'd1);

assign xor_ln302_152_fu_39754_p2 = (p_Result_394_fu_39722_p3 ^ p_Result_393_fu_39708_p3);

assign xor_ln302_153_fu_39760_p2 = (xor_ln302_152_fu_39754_p2 ^ 1'd1);

assign xor_ln302_154_fu_39856_p2 = (p_Result_396_fu_39824_p3 ^ p_Result_395_fu_39810_p3);

assign xor_ln302_155_fu_39862_p2 = (xor_ln302_154_fu_39856_p2 ^ 1'd1);

assign xor_ln302_156_fu_39958_p2 = (p_Result_398_fu_39926_p3 ^ p_Result_397_fu_39912_p3);

assign xor_ln302_157_fu_39964_p2 = (xor_ln302_156_fu_39958_p2 ^ 1'd1);

assign xor_ln302_158_fu_40060_p2 = (p_Result_400_fu_40028_p3 ^ p_Result_399_fu_40014_p3);

assign xor_ln302_159_fu_40066_p2 = (xor_ln302_158_fu_40060_p2 ^ 1'd1);

assign xor_ln302_15_fu_23286_p2 = (xor_ln302_14_fu_23280_p2 ^ 1'd1);

assign xor_ln302_160_fu_40162_p2 = (p_Result_402_fu_40130_p3 ^ p_Result_401_fu_40116_p3);

assign xor_ln302_161_fu_40168_p2 = (xor_ln302_160_fu_40162_p2 ^ 1'd1);

assign xor_ln302_16_fu_23378_p2 = (p_Result_258_fu_23346_p3 ^ p_Result_257_fu_23332_p3);

assign xor_ln302_17_fu_23384_p2 = (xor_ln302_16_fu_23378_p2 ^ 1'd1);

assign xor_ln302_18_fu_23480_p2 = (p_Result_260_fu_23448_p3 ^ p_Result_259_fu_23434_p3);

assign xor_ln302_19_fu_23486_p2 = (xor_ln302_18_fu_23480_p2 ^ 1'd1);

assign xor_ln302_1_fu_22600_p2 = (xor_ln302_fu_22594_p2 ^ 1'd1);

assign xor_ln302_20_fu_23582_p2 = (p_Result_262_fu_23550_p3 ^ p_Result_261_fu_23536_p3);

assign xor_ln302_21_fu_23588_p2 = (xor_ln302_20_fu_23582_p2 ^ 1'd1);

assign xor_ln302_22_fu_23684_p2 = (p_Result_264_fu_23652_p3 ^ p_Result_263_fu_23638_p3);

assign xor_ln302_23_fu_23690_p2 = (xor_ln302_22_fu_23684_p2 ^ 1'd1);

assign xor_ln302_24_fu_23786_p2 = (p_Result_266_fu_23754_p3 ^ p_Result_265_fu_23740_p3);

assign xor_ln302_25_fu_23792_p2 = (xor_ln302_24_fu_23786_p2 ^ 1'd1);

assign xor_ln302_26_fu_23888_p2 = (p_Result_268_fu_23856_p3 ^ p_Result_267_fu_23842_p3);

assign xor_ln302_27_fu_23894_p2 = (xor_ln302_26_fu_23888_p2 ^ 1'd1);

assign xor_ln302_28_fu_23990_p2 = (p_Result_270_fu_23958_p3 ^ p_Result_269_fu_23944_p3);

assign xor_ln302_29_fu_23996_p2 = (xor_ln302_28_fu_23990_p2 ^ 1'd1);

assign xor_ln302_2_fu_22692_p2 = (p_Result_244_fu_22660_p3 ^ p_Result_243_fu_22646_p3);

assign xor_ln302_30_fu_24092_p2 = (p_Result_272_fu_24060_p3 ^ p_Result_271_fu_24046_p3);

assign xor_ln302_31_fu_24098_p2 = (xor_ln302_30_fu_24092_p2 ^ 1'd1);

assign xor_ln302_32_fu_24194_p2 = (p_Result_274_fu_24162_p3 ^ p_Result_273_fu_24148_p3);

assign xor_ln302_33_fu_24200_p2 = (xor_ln302_32_fu_24194_p2 ^ 1'd1);

assign xor_ln302_34_fu_24296_p2 = (p_Result_276_fu_24264_p3 ^ p_Result_275_fu_24250_p3);

assign xor_ln302_35_fu_24302_p2 = (xor_ln302_34_fu_24296_p2 ^ 1'd1);

assign xor_ln302_36_fu_28481_p2 = (p_Result_278_fu_28449_p3 ^ p_Result_277_fu_28436_p3);

assign xor_ln302_37_fu_28487_p2 = (xor_ln302_36_fu_28481_p2 ^ 1'd1);

assign xor_ln302_38_fu_28581_p2 = (p_Result_280_fu_28549_p3 ^ p_Result_279_fu_28536_p3);

assign xor_ln302_39_fu_28587_p2 = (xor_ln302_38_fu_28581_p2 ^ 1'd1);

assign xor_ln302_3_fu_22698_p2 = (xor_ln302_2_fu_22692_p2 ^ 1'd1);

assign xor_ln302_40_fu_28643_p2 = (p_Result_282_reg_41729 ^ p_Result_281_reg_41716);

assign xor_ln302_41_fu_28647_p2 = (xor_ln302_40_fu_28643_p2 ^ 1'd1);

assign xor_ln302_42_fu_28739_p2 = (p_Result_284_fu_28707_p3 ^ p_Result_283_fu_28694_p3);

assign xor_ln302_43_fu_28745_p2 = (xor_ln302_42_fu_28739_p2 ^ 1'd1);

assign xor_ln302_44_fu_28839_p2 = (p_Result_286_fu_28807_p3 ^ p_Result_285_fu_28794_p3);

assign xor_ln302_45_fu_28845_p2 = (xor_ln302_44_fu_28839_p2 ^ 1'd1);

assign xor_ln302_46_fu_28939_p2 = (p_Result_288_fu_28907_p3 ^ p_Result_287_fu_28894_p3);

assign xor_ln302_47_fu_28945_p2 = (xor_ln302_46_fu_28939_p2 ^ 1'd1);

assign xor_ln302_48_fu_29001_p2 = (p_Result_290_reg_41749 ^ p_Result_289_reg_41736);

assign xor_ln302_49_fu_29005_p2 = (xor_ln302_48_fu_29001_p2 ^ 1'd1);

assign xor_ln302_4_fu_22790_p2 = (p_Result_246_fu_22758_p3 ^ p_Result_245_fu_22744_p3);

assign xor_ln302_50_fu_29097_p2 = (p_Result_292_fu_29065_p3 ^ p_Result_291_fu_29052_p3);

assign xor_ln302_51_fu_29103_p2 = (xor_ln302_50_fu_29097_p2 ^ 1'd1);

assign xor_ln302_52_fu_29197_p2 = (p_Result_294_fu_29165_p3 ^ p_Result_293_fu_29152_p3);

assign xor_ln302_53_fu_29203_p2 = (xor_ln302_52_fu_29197_p2 ^ 1'd1);

assign xor_ln302_54_fu_29299_p2 = (p_Result_296_fu_29267_p3 ^ p_Result_295_fu_29253_p3);

assign xor_ln302_55_fu_29305_p2 = (xor_ln302_54_fu_29299_p2 ^ 1'd1);

assign xor_ln302_56_fu_29401_p2 = (p_Result_298_fu_29369_p3 ^ p_Result_297_fu_29355_p3);

assign xor_ln302_57_fu_29407_p2 = (xor_ln302_56_fu_29401_p2 ^ 1'd1);

assign xor_ln302_58_fu_29503_p2 = (p_Result_300_fu_29471_p3 ^ p_Result_299_fu_29457_p3);

assign xor_ln302_59_fu_29509_p2 = (xor_ln302_58_fu_29503_p2 ^ 1'd1);

assign xor_ln302_5_fu_22796_p2 = (xor_ln302_4_fu_22790_p2 ^ 1'd1);

assign xor_ln302_60_fu_29605_p2 = (p_Result_302_fu_29573_p3 ^ p_Result_301_fu_29559_p3);

assign xor_ln302_61_fu_29611_p2 = (xor_ln302_60_fu_29605_p2 ^ 1'd1);

assign xor_ln302_62_fu_29707_p2 = (p_Result_304_fu_29675_p3 ^ p_Result_303_fu_29661_p3);

assign xor_ln302_63_fu_29713_p2 = (xor_ln302_62_fu_29707_p2 ^ 1'd1);

assign xor_ln302_64_fu_29809_p2 = (p_Result_306_fu_29777_p3 ^ p_Result_305_fu_29763_p3);

assign xor_ln302_65_fu_29815_p2 = (xor_ln302_64_fu_29809_p2 ^ 1'd1);

assign xor_ln302_66_fu_29911_p2 = (p_Result_308_fu_29879_p3 ^ p_Result_307_fu_29865_p3);

assign xor_ln302_67_fu_29917_p2 = (xor_ln302_66_fu_29911_p2 ^ 1'd1);

assign xor_ln302_68_fu_30013_p2 = (p_Result_310_fu_29981_p3 ^ p_Result_309_fu_29967_p3);

assign xor_ln302_69_fu_30019_p2 = (xor_ln302_68_fu_30013_p2 ^ 1'd1);

assign xor_ln302_6_fu_22888_p2 = (p_Result_248_fu_22856_p3 ^ p_Result_247_fu_22842_p3);

assign xor_ln302_70_fu_30115_p2 = (p_Result_312_fu_30083_p3 ^ p_Result_311_fu_30069_p3);

assign xor_ln302_71_fu_30121_p2 = (xor_ln302_70_fu_30115_p2 ^ 1'd1);

assign xor_ln302_72_fu_33942_p2 = (p_Result_314_reg_42247 ^ p_Result_313_reg_42234);

assign xor_ln302_73_fu_33946_p2 = (xor_ln302_72_fu_33942_p2 ^ 1'd1);

assign xor_ln302_74_fu_34000_p2 = (p_Result_316_reg_42267 ^ p_Result_315_reg_42254);

assign xor_ln302_75_fu_34004_p2 = (xor_ln302_74_fu_34000_p2 ^ 1'd1);

assign xor_ln302_76_fu_30289_p2 = (p_Result_318_fu_30257_p3 ^ p_Result_317_fu_30243_p3);

assign xor_ln302_77_fu_30295_p2 = (xor_ln302_76_fu_30289_p2 ^ 1'd1);

assign xor_ln302_78_fu_34058_p2 = (p_Result_320_reg_42293 ^ p_Result_319_reg_42280);

assign xor_ln302_79_fu_34062_p2 = (xor_ln302_78_fu_34058_p2 ^ 1'd1);

assign xor_ln302_7_fu_22894_p2 = (xor_ln302_6_fu_22888_p2 ^ 1'd1);

assign xor_ln302_80_fu_34116_p2 = (p_Result_322_reg_42313 ^ p_Result_321_reg_42300);

assign xor_ln302_81_fu_34120_p2 = (xor_ln302_80_fu_34116_p2 ^ 1'd1);

assign xor_ln302_82_fu_34174_p2 = (p_Result_324_reg_42333 ^ p_Result_323_reg_42320);

assign xor_ln302_83_fu_34178_p2 = (xor_ln302_82_fu_34174_p2 ^ 1'd1);

assign xor_ln302_84_fu_30499_p2 = (p_Result_326_fu_30467_p3 ^ p_Result_325_fu_30453_p3);

assign xor_ln302_85_fu_30505_p2 = (xor_ln302_84_fu_30499_p2 ^ 1'd1);

assign xor_ln302_86_fu_34232_p2 = (p_Result_328_reg_42359 ^ p_Result_327_reg_42346);

assign xor_ln302_87_fu_34236_p2 = (xor_ln302_86_fu_34232_p2 ^ 1'd1);

assign xor_ln302_88_fu_34290_p2 = (p_Result_330_reg_42379 ^ p_Result_329_reg_42366);

assign xor_ln302_89_fu_34294_p2 = (xor_ln302_88_fu_34290_p2 ^ 1'd1);

assign xor_ln302_8_fu_22986_p2 = (p_Result_250_fu_22954_p3 ^ p_Result_249_fu_22940_p3);

assign xor_ln302_90_fu_34388_p2 = (p_Result_332_fu_34356_p3 ^ p_Result_331_fu_34342_p3);

assign xor_ln302_91_fu_34394_p2 = (xor_ln302_90_fu_34388_p2 ^ 1'd1);

assign xor_ln302_92_fu_34490_p2 = (p_Result_334_fu_34458_p3 ^ p_Result_333_fu_34444_p3);

assign xor_ln302_93_fu_34496_p2 = (xor_ln302_92_fu_34490_p2 ^ 1'd1);

assign xor_ln302_94_fu_34590_p2 = (p_Result_336_fu_34558_p3 ^ p_Result_335_fu_34545_p3);

assign xor_ln302_95_fu_34596_p2 = (xor_ln302_94_fu_34590_p2 ^ 1'd1);

assign xor_ln302_96_fu_34692_p2 = (p_Result_338_fu_34660_p3 ^ p_Result_337_fu_34646_p3);

assign xor_ln302_97_fu_34698_p2 = (xor_ln302_96_fu_34692_p2 ^ 1'd1);

assign xor_ln302_98_fu_34794_p2 = (p_Result_340_fu_34762_p3 ^ p_Result_339_fu_34748_p3);

assign xor_ln302_99_fu_34800_p2 = (xor_ln302_98_fu_34794_p2 ^ 1'd1);

assign xor_ln302_9_fu_22992_p2 = (xor_ln302_8_fu_22986_p2 ^ 1'd1);

assign xor_ln302_fu_22594_p2 = (p_Result_242_fu_22562_p3 ^ p_Result_241_fu_22548_p3);

assign xor_ln888_101_fu_31285_p2 = (p_Result_155_reg_41947 ^ 1'd1);

assign xor_ln888_103_fu_27755_p2 = (p_Result_158_fu_27701_p3 ^ 1'd1);

assign xor_ln888_105_fu_31449_p2 = (p_Result_161_reg_41998 ^ 1'd1);

assign xor_ln888_107_fu_31598_p2 = (p_Result_164_reg_42027 ^ 1'd1);

assign xor_ln888_109_fu_31747_p2 = (p_Result_167_reg_42056 ^ 1'd1);

assign xor_ln888_111_fu_31896_p2 = (p_Result_170_reg_42085 ^ 1'd1);

assign xor_ln888_113_fu_32045_p2 = (p_Result_173_reg_42114 ^ 1'd1);

assign xor_ln888_115_fu_32194_p2 = (p_Result_176_reg_42143 ^ 1'd1);

assign xor_ln888_117_fu_32343_p2 = (p_Result_179_reg_42172 ^ 1'd1);

assign xor_ln888_119_fu_28277_p2 = (p_Result_182_fu_28223_p3 ^ 1'd1);

assign xor_ln888_11_fu_18894_p2 = (p_Result_13_reg_40437 ^ 1'd1);

assign xor_ln888_121_fu_32509_p2 = (p_Result_185_reg_42216 ^ 1'd1);

assign xor_ln888_123_fu_36173_p2 = (p_Result_188_reg_42392 ^ 1'd1);

assign xor_ln888_125_fu_36298_p2 = (p_Result_191_reg_42423 ^ 1'd1);

assign xor_ln888_127_fu_36423_p2 = (p_Result_194_reg_42454 ^ 1'd1);

assign xor_ln888_129_fu_36548_p2 = (p_Result_197_reg_42485 ^ 1'd1);

assign xor_ln888_131_fu_36673_p2 = (p_Result_200_reg_42516 ^ 1'd1);

assign xor_ln888_133_fu_33053_p2 = (p_Result_203_fu_32999_p3 ^ 1'd1);

assign xor_ln888_135_fu_36815_p2 = (p_Result_206_reg_42562 ^ 1'd1);

assign xor_ln888_137_fu_36940_p2 = (p_Result_209_reg_42593 ^ 1'd1);

assign xor_ln888_139_fu_37065_p2 = (p_Result_212_reg_42624 ^ 1'd1);

assign xor_ln888_13_fu_19019_p2 = (p_Result_16_reg_40468 ^ 1'd1);

assign xor_ln888_141_fu_37212_p2 = (p_Result_215_reg_42660 ^ 1'd1);

assign xor_ln888_143_fu_37361_p2 = (p_Result_218_reg_42689 ^ 1'd1);

assign xor_ln888_145_fu_37510_p2 = (p_Result_221_reg_42718 ^ 1'd1);

assign xor_ln888_147_fu_37659_p2 = (p_Result_224_reg_42747 ^ 1'd1);

assign xor_ln888_149_fu_33650_p2 = (p_Result_227_fu_33596_p3 ^ 1'd1);

assign xor_ln888_151_fu_37825_p2 = (p_Result_230_reg_42791 ^ 1'd1);

assign xor_ln888_153_fu_37974_p2 = (p_Result_233_reg_42820 ^ 1'd1);

assign xor_ln888_155_fu_38123_p2 = (p_Result_236_reg_42849 ^ 1'd1);

assign xor_ln888_157_fu_38272_p2 = (p_Result_239_reg_42878 ^ 1'd1);

assign xor_ln888_15_fu_16901_p2 = (p_Result_19_fu_16847_p3 ^ 1'd1);

assign xor_ln888_17_fu_19158_p2 = (p_Result_22_reg_40514 ^ 1'd1);

assign xor_ln888_19_fu_19282_p2 = (p_Result_25_reg_40545 ^ 1'd1);

assign xor_ln888_1_fu_18502_p2 = (p_Result_1_reg_40329 ^ 1'd1);

assign xor_ln888_21_fu_19429_p2 = (p_Result_28_reg_40581 ^ 1'd1);

assign xor_ln888_23_fu_19612_p2 = (p_Result_36_reg_40640 ^ 1'd1);

assign xor_ln888_25_fu_19761_p2 = (p_Result_39_reg_40669 ^ 1'd1);

assign xor_ln888_27_fu_19905_p2 = (p_Result_44_reg_40708 ^ 1'd1);

assign xor_ln888_29_fu_20052_p2 = (p_Result_47_reg_40744 ^ 1'd1);

assign xor_ln888_2_fu_17423_p2 = (p_Result_33_fu_17383_p3 ^ 1'd1);

assign xor_ln888_31_fu_20201_p2 = (p_Result_50_reg_40773 ^ 1'd1);

assign xor_ln888_33_fu_20346_p2 = (p_Result_53_reg_40802 ^ 1'd1);

assign xor_ln888_35_fu_20475_p2 = (p_Result_56_reg_40831 ^ 1'd1);

assign xor_ln888_37_fu_20608_p2 = (p_Result_59_reg_40860 ^ 1'd1);

assign xor_ln888_39_fu_20753_p2 = (p_Result_62_reg_40889 ^ 1'd1);

assign xor_ln888_41_fu_20882_p2 = (p_Result_65_reg_40918 ^ 1'd1);

assign xor_ln888_43_fu_21011_p2 = (p_Result_68_reg_40947 ^ 1'd1);

assign xor_ln888_45_fu_18275_p2 = (p_Result_71_fu_18221_p3 ^ 1'd1);

assign xor_ln888_47_fu_21157_p2 = (p_Result_74_reg_40991 ^ 1'd1);

assign xor_ln888_49_fu_21286_p2 = (p_Result_77_reg_41020 ^ 1'd1);

assign xor_ln888_4_fu_17651_p2 = (p_Result_41_fu_17611_p3 ^ 1'd1);

assign xor_ln888_51_fu_24539_p2 = (p_Result_80_reg_41154 ^ 1'd1);

assign xor_ln888_53_fu_24663_p2 = (p_Result_83_reg_41185 ^ 1'd1);

assign xor_ln888_55_fu_24788_p2 = (p_Result_86_reg_41216 ^ 1'd1);

assign xor_ln888_57_fu_24913_p2 = (p_Result_89_reg_41247 ^ 1'd1);

assign xor_ln888_59_fu_25038_p2 = (p_Result_92_reg_41278 ^ 1'd1);

assign xor_ln888_5_fu_18627_p2 = (p_Result_4_reg_40360 ^ 1'd1);

assign xor_ln888_61_fu_25163_p2 = (p_Result_95_reg_41309 ^ 1'd1);

assign xor_ln888_63_fu_25288_p2 = (p_Result_98_reg_41340 ^ 1'd1);

assign xor_ln888_65_fu_25413_p2 = (p_Result_101_reg_41371 ^ 1'd1);

assign xor_ln888_67_fu_25535_p2 = (p_Result_104_reg_41402 ^ 1'd1);

assign xor_ln888_69_fu_25681_p2 = (p_Result_107_reg_41438 ^ 1'd1);

assign xor_ln888_71_fu_25830_p2 = (p_Result_110_reg_41467 ^ 1'd1);

assign xor_ln888_73_fu_25979_p2 = (p_Result_113_reg_41496 ^ 1'd1);

assign xor_ln888_75_fu_22224_p2 = (p_Result_116_fu_22170_p3 ^ 1'd1);

assign xor_ln888_77_fu_26145_p2 = (p_Result_119_reg_41540 ^ 1'd1);

assign xor_ln888_79_fu_26294_p2 = (p_Result_122_reg_41569 ^ 1'd1);

assign xor_ln888_7_fu_16523_p2 = (p_Result_7_fu_16469_p3 ^ 1'd1);

assign xor_ln888_81_fu_26443_p2 = (p_Result_125_reg_41598 ^ 1'd1);

assign xor_ln888_83_fu_26592_p2 = (p_Result_128_reg_41627 ^ 1'd1);

assign xor_ln888_85_fu_26741_p2 = (p_Result_131_reg_41656 ^ 1'd1);

assign xor_ln888_87_fu_26960_p2 = (p_Result_134_fu_26915_p3 ^ 1'd1);

assign xor_ln888_89_fu_30643_p2 = (p_Result_137_reg_41777 ^ 1'd1);

assign xor_ln888_91_fu_30768_p2 = (p_Result_140_reg_41808 ^ 1'd1);

assign xor_ln888_93_fu_30893_p2 = (p_Result_143_reg_41839 ^ 1'd1);

assign xor_ln888_95_fu_31018_p2 = (p_Result_146_reg_41870 ^ 1'd1);

assign xor_ln888_97_fu_31143_p2 = (p_Result_149_reg_41901 ^ 1'd1);

assign xor_ln888_99_fu_27494_p2 = (p_Result_152_fu_27440_p3 ^ 1'd1);

assign xor_ln888_9_fu_18769_p2 = (p_Result_10_reg_40406 ^ 1'd1);

assign xor_ln888_fu_17259_p2 = (p_Result_31_fu_17211_p3 ^ 1'd1);

assign xor_ln890_10_fu_17279_p2 = (tmp_63_fu_17271_p3 ^ 1'd1);

assign xor_ln890_11_fu_19636_p2 = (tmp_72_fu_19628_p3 ^ 1'd1);

assign xor_ln890_12_fu_19785_p2 = (tmp_78_fu_19777_p3 ^ 1'd1);

assign xor_ln890_13_fu_19928_p2 = (tmp_87_fu_19920_p3 ^ 1'd1);

assign xor_ln890_14_fu_20076_p2 = (tmp_93_fu_20068_p3 ^ 1'd1);

assign xor_ln890_15_fu_20225_p2 = (tmp_99_fu_20217_p3 ^ 1'd1);

assign xor_ln890_16_fu_20370_p2 = (tmp_105_fu_20362_p3 ^ 1'd1);

assign xor_ln890_17_fu_20499_p2 = (tmp_111_fu_20491_p3 ^ 1'd1);

assign xor_ln890_18_fu_20632_p2 = (tmp_117_fu_20624_p3 ^ 1'd1);

assign xor_ln890_19_fu_20777_p2 = (tmp_123_fu_20769_p3 ^ 1'd1);

assign xor_ln890_1_fu_18650_p2 = (tmp_9_fu_18642_p3 ^ 1'd1);

assign xor_ln890_20_fu_20906_p2 = (tmp_129_fu_20898_p3 ^ 1'd1);

assign xor_ln890_21_fu_21035_p2 = (tmp_135_fu_21027_p3 ^ 1'd1);

assign xor_ln890_22_fu_18301_p2 = (tmp_141_fu_18293_p3 ^ 1'd1);

assign xor_ln890_23_fu_21181_p2 = (tmp_147_fu_21173_p3 ^ 1'd1);

assign xor_ln890_24_fu_21310_p2 = (tmp_153_fu_21302_p3 ^ 1'd1);

assign xor_ln890_25_fu_24562_p2 = (tmp_159_fu_24554_p3 ^ 1'd1);

assign xor_ln890_26_fu_24686_p2 = (tmp_165_fu_24678_p3 ^ 1'd1);

assign xor_ln890_27_fu_24811_p2 = (tmp_171_fu_24803_p3 ^ 1'd1);

assign xor_ln890_28_fu_24936_p2 = (tmp_177_fu_24928_p3 ^ 1'd1);

assign xor_ln890_29_fu_25061_p2 = (tmp_183_fu_25053_p3 ^ 1'd1);

assign xor_ln890_2_fu_16549_p2 = (tmp_15_fu_16541_p3 ^ 1'd1);

assign xor_ln890_30_fu_25186_p2 = (tmp_189_fu_25178_p3 ^ 1'd1);

assign xor_ln890_31_fu_25311_p2 = (tmp_195_fu_25303_p3 ^ 1'd1);

assign xor_ln890_32_fu_25436_p2 = (tmp_201_fu_25428_p3 ^ 1'd1);

assign xor_ln890_33_fu_25558_p2 = (tmp_207_fu_25550_p3 ^ 1'd1);

assign xor_ln890_34_fu_25705_p2 = (tmp_213_fu_25697_p3 ^ 1'd1);

assign xor_ln890_35_fu_25854_p2 = (tmp_219_fu_25846_p3 ^ 1'd1);

assign xor_ln890_36_fu_26003_p2 = (tmp_225_fu_25995_p3 ^ 1'd1);

assign xor_ln890_37_fu_22250_p2 = (tmp_231_fu_22242_p3 ^ 1'd1);

assign xor_ln890_38_fu_26169_p2 = (tmp_237_fu_26161_p3 ^ 1'd1);

assign xor_ln890_39_fu_26318_p2 = (tmp_243_fu_26310_p3 ^ 1'd1);

assign xor_ln890_3_fu_18792_p2 = (tmp_21_fu_18784_p3 ^ 1'd1);

assign xor_ln890_40_fu_26467_p2 = (tmp_249_fu_26459_p3 ^ 1'd1);

assign xor_ln890_41_fu_26616_p2 = (tmp_255_fu_26608_p3 ^ 1'd1);

assign xor_ln890_42_fu_26765_p2 = (tmp_261_fu_26757_p3 ^ 1'd1);

assign xor_ln890_43_fu_26986_p2 = (tmp_267_fu_26978_p3 ^ 1'd1);

assign xor_ln890_44_fu_30666_p2 = (tmp_273_fu_30658_p3 ^ 1'd1);

assign xor_ln890_45_fu_30791_p2 = (tmp_279_fu_30783_p3 ^ 1'd1);

assign xor_ln890_46_fu_30916_p2 = (tmp_285_fu_30908_p3 ^ 1'd1);

assign xor_ln890_47_fu_31041_p2 = (tmp_291_fu_31033_p3 ^ 1'd1);

assign xor_ln890_48_fu_31166_p2 = (tmp_297_fu_31158_p3 ^ 1'd1);

assign xor_ln890_49_fu_27520_p2 = (tmp_303_fu_27512_p3 ^ 1'd1);

assign xor_ln890_4_fu_18917_p2 = (tmp_27_fu_18909_p3 ^ 1'd1);

assign xor_ln890_50_fu_31308_p2 = (tmp_309_fu_31300_p3 ^ 1'd1);

assign xor_ln890_51_fu_27781_p2 = (tmp_315_fu_27773_p3 ^ 1'd1);

assign xor_ln890_52_fu_31473_p2 = (tmp_321_fu_31465_p3 ^ 1'd1);

assign xor_ln890_53_fu_31622_p2 = (tmp_327_fu_31614_p3 ^ 1'd1);

assign xor_ln890_54_fu_31771_p2 = (tmp_333_fu_31763_p3 ^ 1'd1);

assign xor_ln890_55_fu_31920_p2 = (tmp_339_fu_31912_p3 ^ 1'd1);

assign xor_ln890_56_fu_32069_p2 = (tmp_345_fu_32061_p3 ^ 1'd1);

assign xor_ln890_57_fu_32218_p2 = (tmp_351_fu_32210_p3 ^ 1'd1);

assign xor_ln890_58_fu_32367_p2 = (tmp_357_fu_32359_p3 ^ 1'd1);

assign xor_ln890_59_fu_28303_p2 = (tmp_363_fu_28295_p3 ^ 1'd1);

assign xor_ln890_5_fu_19042_p2 = (tmp_33_fu_19034_p3 ^ 1'd1);

assign xor_ln890_60_fu_32533_p2 = (tmp_369_fu_32525_p3 ^ 1'd1);

assign xor_ln890_61_fu_36196_p2 = (tmp_375_fu_36188_p3 ^ 1'd1);

assign xor_ln890_62_fu_36321_p2 = (tmp_381_fu_36313_p3 ^ 1'd1);

assign xor_ln890_63_fu_36446_p2 = (tmp_387_fu_36438_p3 ^ 1'd1);

assign xor_ln890_64_fu_36571_p2 = (tmp_393_fu_36563_p3 ^ 1'd1);

assign xor_ln890_65_fu_36696_p2 = (tmp_399_fu_36688_p3 ^ 1'd1);

assign xor_ln890_66_fu_33079_p2 = (tmp_405_fu_33071_p3 ^ 1'd1);

assign xor_ln890_67_fu_36838_p2 = (tmp_411_fu_36830_p3 ^ 1'd1);

assign xor_ln890_68_fu_36963_p2 = (tmp_417_fu_36955_p3 ^ 1'd1);

assign xor_ln890_69_fu_37088_p2 = (tmp_423_fu_37080_p3 ^ 1'd1);

assign xor_ln890_6_fu_16927_p2 = (tmp_39_fu_16919_p3 ^ 1'd1);

assign xor_ln890_70_fu_37236_p2 = (tmp_429_fu_37228_p3 ^ 1'd1);

assign xor_ln890_71_fu_37385_p2 = (tmp_435_fu_37377_p3 ^ 1'd1);

assign xor_ln890_72_fu_37534_p2 = (tmp_441_fu_37526_p3 ^ 1'd1);

assign xor_ln890_73_fu_37683_p2 = (tmp_447_fu_37675_p3 ^ 1'd1);

assign xor_ln890_74_fu_33676_p2 = (tmp_453_fu_33668_p3 ^ 1'd1);

assign xor_ln890_75_fu_37849_p2 = (tmp_459_fu_37841_p3 ^ 1'd1);

assign xor_ln890_76_fu_37998_p2 = (tmp_465_fu_37990_p3 ^ 1'd1);

assign xor_ln890_77_fu_38147_p2 = (tmp_471_fu_38139_p3 ^ 1'd1);

assign xor_ln890_78_fu_38296_p2 = (tmp_477_fu_38288_p3 ^ 1'd1);

assign xor_ln890_7_fu_19181_p2 = (tmp_45_fu_19173_p3 ^ 1'd1);

assign xor_ln890_8_fu_19305_p2 = (tmp_51_fu_19297_p3 ^ 1'd1);

assign xor_ln890_9_fu_19453_p2 = (tmp_57_fu_19445_p3 ^ 1'd1);

assign xor_ln890_fu_18525_p2 = (tmp_3_fu_18517_p3 ^ 1'd1);

assign xor_ln895_100_fu_31188_p2 = (deleted_zeros_47_fu_31153_p2 ^ 1'd1);

assign xor_ln895_101_fu_31199_p2 = (p_Result_148_reg_41895 ^ 1'd1);

assign xor_ln895_102_fu_27544_p2 = (deleted_zeros_48_fu_27506_p2 ^ 1'd1);

assign xor_ln895_103_fu_27556_p2 = (p_Result_151_fu_27418_p3 ^ 1'd1);

assign xor_ln895_104_fu_31330_p2 = (deleted_zeros_49_fu_31295_p2 ^ 1'd1);

assign xor_ln895_105_fu_31341_p2 = (p_Result_154_reg_41941 ^ 1'd1);

assign xor_ln895_106_fu_27805_p2 = (deleted_zeros_50_fu_27767_p2 ^ 1'd1);

assign xor_ln895_107_fu_27817_p2 = (p_Result_157_fu_27679_p3 ^ 1'd1);

assign xor_ln895_108_fu_31495_p2 = (deleted_zeros_51_fu_31460_p2 ^ 1'd1);

assign xor_ln895_109_fu_31507_p2 = (p_Result_160_reg_41987 ^ 1'd1);

assign xor_ln895_10_fu_19064_p2 = (deleted_zeros_5_fu_19029_p2 ^ 1'd1);

assign xor_ln895_110_fu_31644_p2 = (deleted_zeros_52_fu_31609_p2 ^ 1'd1);

assign xor_ln895_111_fu_31656_p2 = (p_Result_163_reg_42016 ^ 1'd1);

assign xor_ln895_112_fu_31793_p2 = (deleted_zeros_53_fu_31758_p2 ^ 1'd1);

assign xor_ln895_113_fu_31805_p2 = (p_Result_166_reg_42045 ^ 1'd1);

assign xor_ln895_114_fu_31942_p2 = (deleted_zeros_54_fu_31907_p2 ^ 1'd1);

assign xor_ln895_115_fu_31954_p2 = (p_Result_169_reg_42074 ^ 1'd1);

assign xor_ln895_116_fu_32091_p2 = (deleted_zeros_55_fu_32056_p2 ^ 1'd1);

assign xor_ln895_117_fu_32103_p2 = (p_Result_172_reg_42103 ^ 1'd1);

assign xor_ln895_118_fu_32240_p2 = (deleted_zeros_56_fu_32205_p2 ^ 1'd1);

assign xor_ln895_119_fu_32252_p2 = (p_Result_175_reg_42132 ^ 1'd1);

assign xor_ln895_11_fu_19075_p2 = (p_Result_15_reg_40462 ^ 1'd1);

assign xor_ln895_120_fu_32389_p2 = (deleted_zeros_57_fu_32354_p2 ^ 1'd1);

assign xor_ln895_121_fu_32401_p2 = (p_Result_178_reg_42161 ^ 1'd1);

assign xor_ln895_122_fu_28327_p2 = (deleted_zeros_58_fu_28289_p2 ^ 1'd1);

assign xor_ln895_123_fu_28339_p2 = (p_Result_181_fu_28201_p3 ^ 1'd1);

assign xor_ln895_124_fu_32555_p2 = (deleted_zeros_59_fu_32520_p2 ^ 1'd1);

assign xor_ln895_125_fu_32567_p2 = (p_Result_184_reg_42205 ^ 1'd1);

assign xor_ln895_126_fu_36218_p2 = (deleted_zeros_60_fu_36183_p2 ^ 1'd1);

assign xor_ln895_127_fu_36229_p2 = (p_Result_187_reg_42386 ^ 1'd1);

assign xor_ln895_128_fu_36343_p2 = (deleted_zeros_61_fu_36308_p2 ^ 1'd1);

assign xor_ln895_129_fu_36354_p2 = (p_Result_190_reg_42417 ^ 1'd1);

assign xor_ln895_12_fu_16951_p2 = (deleted_zeros_6_fu_16913_p2 ^ 1'd1);

assign xor_ln895_130_fu_36468_p2 = (deleted_zeros_62_fu_36433_p2 ^ 1'd1);

assign xor_ln895_131_fu_36479_p2 = (p_Result_193_reg_42448 ^ 1'd1);

assign xor_ln895_132_fu_36593_p2 = (deleted_zeros_63_fu_36558_p2 ^ 1'd1);

assign xor_ln895_133_fu_36604_p2 = (p_Result_196_reg_42479 ^ 1'd1);

assign xor_ln895_134_fu_36718_p2 = (deleted_zeros_64_fu_36683_p2 ^ 1'd1);

assign xor_ln895_135_fu_36729_p2 = (p_Result_199_reg_42510 ^ 1'd1);

assign xor_ln895_136_fu_33103_p2 = (deleted_zeros_65_fu_33065_p2 ^ 1'd1);

assign xor_ln895_137_fu_33115_p2 = (p_Result_202_fu_32977_p3 ^ 1'd1);

assign xor_ln895_138_fu_36860_p2 = (deleted_zeros_66_fu_36825_p2 ^ 1'd1);

assign xor_ln895_139_fu_36871_p2 = (p_Result_205_reg_42556 ^ 1'd1);

assign xor_ln895_13_fu_16963_p2 = (p_Result_18_fu_16825_p3 ^ 1'd1);

assign xor_ln895_140_fu_36985_p2 = (deleted_zeros_67_fu_36950_p2 ^ 1'd1);

assign xor_ln895_141_fu_36996_p2 = (p_Result_208_reg_42587 ^ 1'd1);

assign xor_ln895_142_fu_37110_p2 = (deleted_zeros_68_fu_37075_p2 ^ 1'd1);

assign xor_ln895_143_fu_37121_p2 = (p_Result_211_reg_42618 ^ 1'd1);

assign xor_ln895_144_fu_37258_p2 = (deleted_zeros_69_fu_37223_p2 ^ 1'd1);

assign xor_ln895_145_fu_37270_p2 = (p_Result_214_reg_42649 ^ 1'd1);

assign xor_ln895_146_fu_37407_p2 = (deleted_zeros_70_fu_37372_p2 ^ 1'd1);

assign xor_ln895_147_fu_37419_p2 = (p_Result_217_reg_42678 ^ 1'd1);

assign xor_ln895_148_fu_37556_p2 = (deleted_zeros_71_fu_37521_p2 ^ 1'd1);

assign xor_ln895_149_fu_37568_p2 = (p_Result_220_reg_42707 ^ 1'd1);

assign xor_ln895_14_fu_19203_p2 = (deleted_zeros_7_fu_19168_p2 ^ 1'd1);

assign xor_ln895_150_fu_37705_p2 = (deleted_zeros_72_fu_37670_p2 ^ 1'd1);

assign xor_ln895_151_fu_37717_p2 = (p_Result_223_reg_42736 ^ 1'd1);

assign xor_ln895_152_fu_33700_p2 = (deleted_zeros_73_fu_33662_p2 ^ 1'd1);

assign xor_ln895_153_fu_33712_p2 = (p_Result_226_fu_33574_p3 ^ 1'd1);

assign xor_ln895_154_fu_37871_p2 = (deleted_zeros_74_fu_37836_p2 ^ 1'd1);

assign xor_ln895_155_fu_37883_p2 = (p_Result_229_reg_42780 ^ 1'd1);

assign xor_ln895_156_fu_38020_p2 = (deleted_zeros_75_fu_37985_p2 ^ 1'd1);

assign xor_ln895_157_fu_38032_p2 = (p_Result_232_reg_42809 ^ 1'd1);

assign xor_ln895_158_fu_38169_p2 = (deleted_zeros_76_fu_38134_p2 ^ 1'd1);

assign xor_ln895_159_fu_38181_p2 = (p_Result_235_reg_42838 ^ 1'd1);

assign xor_ln895_15_fu_19214_p2 = (p_Result_21_reg_40508 ^ 1'd1);

assign xor_ln895_160_fu_38318_p2 = (deleted_zeros_77_fu_38283_p2 ^ 1'd1);

assign xor_ln895_161_fu_38330_p2 = (p_Result_238_reg_42867 ^ 1'd1);

assign xor_ln895_162_fu_22570_p2 = (p_Result_241_fu_22548_p3 ^ 1'd1);

assign xor_ln895_163_fu_22668_p2 = (p_Result_243_fu_22646_p3 ^ 1'd1);

assign xor_ln895_164_fu_22766_p2 = (p_Result_245_fu_22744_p3 ^ 1'd1);

assign xor_ln895_165_fu_22864_p2 = (p_Result_247_fu_22842_p3 ^ 1'd1);

assign xor_ln895_166_fu_22962_p2 = (p_Result_249_fu_22940_p3 ^ 1'd1);

assign xor_ln895_167_fu_23060_p2 = (p_Result_251_fu_23038_p3 ^ 1'd1);

assign xor_ln895_168_fu_23158_p2 = (p_Result_253_fu_23136_p3 ^ 1'd1);

assign xor_ln895_169_fu_23256_p2 = (p_Result_255_fu_23234_p3 ^ 1'd1);

assign xor_ln895_16_fu_19327_p2 = (deleted_zeros_8_fu_19292_p2 ^ 1'd1);

assign xor_ln895_170_fu_23354_p2 = (p_Result_257_fu_23332_p3 ^ 1'd1);

assign xor_ln895_171_fu_23456_p2 = (p_Result_259_fu_23434_p3 ^ 1'd1);

assign xor_ln895_172_fu_23558_p2 = (p_Result_261_fu_23536_p3 ^ 1'd1);

assign xor_ln895_173_fu_23660_p2 = (p_Result_263_fu_23638_p3 ^ 1'd1);

assign xor_ln895_174_fu_23762_p2 = (p_Result_265_fu_23740_p3 ^ 1'd1);

assign xor_ln895_175_fu_23864_p2 = (p_Result_267_fu_23842_p3 ^ 1'd1);

assign xor_ln895_176_fu_23966_p2 = (p_Result_269_fu_23944_p3 ^ 1'd1);

assign xor_ln895_177_fu_24068_p2 = (p_Result_271_fu_24046_p3 ^ 1'd1);

assign xor_ln895_178_fu_24170_p2 = (p_Result_273_fu_24148_p3 ^ 1'd1);

assign xor_ln895_179_fu_24272_p2 = (p_Result_275_fu_24250_p3 ^ 1'd1);

assign xor_ln895_17_fu_19338_p2 = (p_Result_24_reg_40539 ^ 1'd1);

assign xor_ln895_180_fu_28457_p2 = (p_Result_277_fu_28436_p3 ^ 1'd1);

assign xor_ln895_181_fu_28557_p2 = (p_Result_279_fu_28536_p3 ^ 1'd1);

assign xor_ln895_182_fu_28623_p2 = (p_Result_281_reg_41716 ^ 1'd1);

assign xor_ln895_183_fu_28715_p2 = (p_Result_283_fu_28694_p3 ^ 1'd1);

assign xor_ln895_184_fu_28815_p2 = (p_Result_285_fu_28794_p3 ^ 1'd1);

assign xor_ln895_185_fu_28915_p2 = (p_Result_287_fu_28894_p3 ^ 1'd1);

assign xor_ln895_186_fu_28981_p2 = (p_Result_289_reg_41736 ^ 1'd1);

assign xor_ln895_187_fu_29073_p2 = (p_Result_291_fu_29052_p3 ^ 1'd1);

assign xor_ln895_188_fu_29173_p2 = (p_Result_293_fu_29152_p3 ^ 1'd1);

assign xor_ln895_189_fu_29275_p2 = (p_Result_295_fu_29253_p3 ^ 1'd1);

assign xor_ln895_18_fu_19475_p2 = (deleted_zeros_9_fu_19440_p2 ^ 1'd1);

assign xor_ln895_190_fu_29377_p2 = (p_Result_297_fu_29355_p3 ^ 1'd1);

assign xor_ln895_191_fu_29479_p2 = (p_Result_299_fu_29457_p3 ^ 1'd1);

assign xor_ln895_192_fu_29581_p2 = (p_Result_301_fu_29559_p3 ^ 1'd1);

assign xor_ln895_193_fu_29683_p2 = (p_Result_303_fu_29661_p3 ^ 1'd1);

assign xor_ln895_194_fu_29785_p2 = (p_Result_305_fu_29763_p3 ^ 1'd1);

assign xor_ln895_195_fu_29887_p2 = (p_Result_307_fu_29865_p3 ^ 1'd1);

assign xor_ln895_196_fu_29989_p2 = (p_Result_309_fu_29967_p3 ^ 1'd1);

assign xor_ln895_197_fu_30091_p2 = (p_Result_311_fu_30069_p3 ^ 1'd1);

assign xor_ln895_198_fu_33922_p2 = (p_Result_313_reg_42234 ^ 1'd1);

assign xor_ln895_199_fu_33980_p2 = (p_Result_315_reg_42254 ^ 1'd1);

assign xor_ln895_19_fu_19487_p2 = (p_Result_27_reg_40570 ^ 1'd1);

assign xor_ln895_1_fu_18558_p2 = (p_Result_s_reg_40323 ^ 1'd1);

assign xor_ln895_200_fu_30265_p2 = (p_Result_317_fu_30243_p3 ^ 1'd1);

assign xor_ln895_201_fu_34038_p2 = (p_Result_319_reg_42280 ^ 1'd1);

assign xor_ln895_202_fu_34096_p2 = (p_Result_321_reg_42300 ^ 1'd1);

assign xor_ln895_203_fu_34154_p2 = (p_Result_323_reg_42320 ^ 1'd1);

assign xor_ln895_204_fu_30475_p2 = (p_Result_325_fu_30453_p3 ^ 1'd1);

assign xor_ln895_205_fu_34212_p2 = (p_Result_327_reg_42346 ^ 1'd1);

assign xor_ln895_206_fu_34270_p2 = (p_Result_329_reg_42366 ^ 1'd1);

assign xor_ln895_207_fu_34364_p2 = (p_Result_331_fu_34342_p3 ^ 1'd1);

assign xor_ln895_208_fu_34466_p2 = (p_Result_333_fu_34444_p3 ^ 1'd1);

assign xor_ln895_209_fu_34566_p2 = (p_Result_335_fu_34545_p3 ^ 1'd1);

assign xor_ln895_20_fu_17315_p2 = (xor_ln895_23_fu_17309_p2 ^ 1'd1);

assign xor_ln895_210_fu_34668_p2 = (p_Result_337_fu_34646_p3 ^ 1'd1);

assign xor_ln895_211_fu_34770_p2 = (p_Result_339_fu_34748_p3 ^ 1'd1);

assign xor_ln895_212_fu_34872_p2 = (p_Result_341_fu_34850_p3 ^ 1'd1);

assign xor_ln895_213_fu_34972_p2 = (p_Result_343_fu_34951_p3 ^ 1'd1);

assign xor_ln895_214_fu_35074_p2 = (p_Result_345_fu_35052_p3 ^ 1'd1);

assign xor_ln895_215_fu_35176_p2 = (p_Result_347_fu_35154_p3 ^ 1'd1);

assign xor_ln895_216_fu_35278_p2 = (p_Result_349_fu_35256_p3 ^ 1'd1);

assign xor_ln895_217_fu_35380_p2 = (p_Result_351_fu_35358_p3 ^ 1'd1);

assign xor_ln895_218_fu_35482_p2 = (p_Result_353_fu_35460_p3 ^ 1'd1);

assign xor_ln895_219_fu_35584_p2 = (p_Result_355_fu_35562_p3 ^ 1'd1);

assign xor_ln895_21_fu_17327_p2 = (p_Result_30_fu_17189_p3 ^ 1'd1);

assign xor_ln895_220_fu_35686_p2 = (p_Result_357_fu_35664_p3 ^ 1'd1);

assign xor_ln895_221_fu_35788_p2 = (p_Result_359_fu_35766_p3 ^ 1'd1);

assign xor_ln895_222_fu_35890_p2 = (p_Result_361_fu_35868_p3 ^ 1'd1);

assign xor_ln895_223_fu_35992_p2 = (p_Result_363_fu_35970_p3 ^ 1'd1);

assign xor_ln895_224_fu_36094_p2 = (p_Result_365_fu_36072_p3 ^ 1'd1);

assign xor_ln895_225_fu_38420_p2 = (p_Result_367_fu_38399_p3 ^ 1'd1);

assign xor_ln895_226_fu_38520_p2 = (p_Result_369_fu_38499_p3 ^ 1'd1);

assign xor_ln895_227_fu_38620_p2 = (p_Result_371_fu_38599_p3 ^ 1'd1);

assign xor_ln895_228_fu_38720_p2 = (p_Result_373_fu_38699_p3 ^ 1'd1);

assign xor_ln895_229_fu_38820_p2 = (p_Result_375_fu_38799_p3 ^ 1'd1);

assign xor_ln895_22_fu_17465_p2 = (xor_ln895_29_fu_17459_p2 ^ 1'd1);

assign xor_ln895_230_fu_38920_p2 = (p_Result_377_fu_38899_p3 ^ 1'd1);

assign xor_ln895_231_fu_39020_p2 = (p_Result_379_fu_38999_p3 ^ 1'd1);

assign xor_ln895_232_fu_39120_p2 = (p_Result_381_fu_39099_p3 ^ 1'd1);

assign xor_ln895_233_fu_39220_p2 = (p_Result_383_fu_39199_p3 ^ 1'd1);

assign xor_ln895_234_fu_39322_p2 = (p_Result_385_fu_39300_p3 ^ 1'd1);

assign xor_ln895_235_fu_39424_p2 = (p_Result_387_fu_39402_p3 ^ 1'd1);

assign xor_ln895_236_fu_39526_p2 = (p_Result_389_fu_39504_p3 ^ 1'd1);

assign xor_ln895_237_fu_39628_p2 = (p_Result_391_fu_39606_p3 ^ 1'd1);

assign xor_ln895_238_fu_39730_p2 = (p_Result_393_fu_39708_p3 ^ 1'd1);

assign xor_ln895_239_fu_39832_p2 = (p_Result_395_fu_39810_p3 ^ 1'd1);

assign xor_ln895_23_fu_17309_p2 = (or_ln888_fu_17265_p2 ^ Range2_all_ones_10_fu_17251_p3);

assign xor_ln895_240_fu_39934_p2 = (p_Result_397_fu_39912_p3 ^ 1'd1);

assign xor_ln895_241_fu_40036_p2 = (p_Result_399_fu_40014_p3 ^ 1'd1);

assign xor_ln895_242_fu_40138_p2 = (p_Result_401_fu_40116_p3 ^ 1'd1);

assign xor_ln895_243_fu_17687_p2 = (or_ln888_2_fu_17657_p2 ^ Range2_all_ones_10_fu_17251_p3);

assign xor_ln895_24_fu_19658_p2 = (deleted_zeros_10_fu_19623_p2 ^ 1'd1);

assign xor_ln895_25_fu_19670_p2 = (p_Result_35_reg_40629 ^ 1'd1);

assign xor_ln895_26_fu_19807_p2 = (deleted_zeros_11_fu_19772_p2 ^ 1'd1);

assign xor_ln895_27_fu_19819_p2 = (p_Result_38_reg_40658 ^ 1'd1);

assign xor_ln895_28_fu_17693_p2 = (xor_ln895_243_fu_17687_p2 ^ 1'd1);

assign xor_ln895_29_fu_17459_p2 = (or_ln888_1_fu_17429_p2 ^ Range2_all_ones_10_fu_17251_p3);

assign xor_ln895_2_fu_18672_p2 = (deleted_zeros_1_fu_18637_p2 ^ 1'd1);

assign xor_ln895_30_fu_19950_p2 = (deleted_zeros_12_fu_19915_p2 ^ 1'd1);

assign xor_ln895_31_fu_19961_p2 = (p_Result_43_reg_40702 ^ 1'd1);

assign xor_ln895_32_fu_20098_p2 = (deleted_zeros_13_fu_20063_p2 ^ 1'd1);

assign xor_ln895_33_fu_20110_p2 = (p_Result_46_reg_40733 ^ 1'd1);

assign xor_ln895_34_fu_20247_p2 = (deleted_zeros_14_fu_20212_p2 ^ 1'd1);

assign xor_ln895_35_fu_20259_p2 = (p_Result_49_reg_40762 ^ 1'd1);

assign xor_ln895_36_fu_20392_p2 = (deleted_zeros_15_fu_20357_p2 ^ 1'd1);

assign xor_ln895_37_fu_20404_p2 = (p_Result_52_reg_40791 ^ 1'd1);

assign xor_ln895_38_fu_20521_p2 = (deleted_zeros_16_fu_20486_p2 ^ 1'd1);

assign xor_ln895_39_fu_20533_p2 = (p_Result_55_reg_40820 ^ 1'd1);

assign xor_ln895_3_fu_18683_p2 = (p_Result_3_reg_40354 ^ 1'd1);

assign xor_ln895_40_fu_20654_p2 = (deleted_zeros_17_fu_20619_p2 ^ 1'd1);

assign xor_ln895_41_fu_20666_p2 = (p_Result_58_reg_40849 ^ 1'd1);

assign xor_ln895_42_fu_20799_p2 = (deleted_zeros_18_fu_20764_p2 ^ 1'd1);

assign xor_ln895_43_fu_20811_p2 = (p_Result_61_reg_40878 ^ 1'd1);

assign xor_ln895_44_fu_20928_p2 = (deleted_zeros_19_fu_20893_p2 ^ 1'd1);

assign xor_ln895_45_fu_20940_p2 = (p_Result_64_reg_40907 ^ 1'd1);

assign xor_ln895_46_fu_21057_p2 = (deleted_zeros_20_fu_21022_p2 ^ 1'd1);

assign xor_ln895_47_fu_21069_p2 = (p_Result_67_reg_40936 ^ 1'd1);

assign xor_ln895_48_fu_18325_p2 = (deleted_zeros_21_fu_18287_p2 ^ 1'd1);

assign xor_ln895_49_fu_18337_p2 = (p_Result_70_fu_18199_p3 ^ 1'd1);

assign xor_ln895_4_fu_16573_p2 = (deleted_zeros_2_fu_16535_p2 ^ 1'd1);

assign xor_ln895_50_fu_21203_p2 = (deleted_zeros_22_fu_21168_p2 ^ 1'd1);

assign xor_ln895_51_fu_21215_p2 = (p_Result_73_reg_40980 ^ 1'd1);

assign xor_ln895_52_fu_21332_p2 = (deleted_zeros_23_fu_21297_p2 ^ 1'd1);

assign xor_ln895_53_fu_21344_p2 = (p_Result_76_reg_41009 ^ 1'd1);

assign xor_ln895_54_fu_24584_p2 = (deleted_zeros_24_fu_24549_p2 ^ 1'd1);

assign xor_ln895_55_fu_24595_p2 = (p_Result_79_reg_41148 ^ 1'd1);

assign xor_ln895_56_fu_24708_p2 = (deleted_zeros_25_fu_24673_p2 ^ 1'd1);

assign xor_ln895_57_fu_24719_p2 = (p_Result_82_reg_41179 ^ 1'd1);

assign xor_ln895_58_fu_24833_p2 = (deleted_zeros_26_fu_24798_p2 ^ 1'd1);

assign xor_ln895_59_fu_24844_p2 = (p_Result_85_reg_41210 ^ 1'd1);

assign xor_ln895_5_fu_16585_p2 = (p_Result_6_fu_16441_p3 ^ 1'd1);

assign xor_ln895_60_fu_24958_p2 = (deleted_zeros_27_fu_24923_p2 ^ 1'd1);

assign xor_ln895_61_fu_24969_p2 = (p_Result_88_reg_41241 ^ 1'd1);

assign xor_ln895_62_fu_25083_p2 = (deleted_zeros_28_fu_25048_p2 ^ 1'd1);

assign xor_ln895_63_fu_25094_p2 = (p_Result_91_reg_41272 ^ 1'd1);

assign xor_ln895_64_fu_25208_p2 = (deleted_zeros_29_fu_25173_p2 ^ 1'd1);

assign xor_ln895_65_fu_25219_p2 = (p_Result_94_reg_41303 ^ 1'd1);

assign xor_ln895_66_fu_25333_p2 = (deleted_zeros_30_fu_25298_p2 ^ 1'd1);

assign xor_ln895_67_fu_25344_p2 = (p_Result_97_reg_41334 ^ 1'd1);

assign xor_ln895_68_fu_25458_p2 = (deleted_zeros_31_fu_25423_p2 ^ 1'd1);

assign xor_ln895_69_fu_25469_p2 = (p_Result_100_reg_41365 ^ 1'd1);

assign xor_ln895_6_fu_18814_p2 = (deleted_zeros_3_fu_18779_p2 ^ 1'd1);

assign xor_ln895_70_fu_25580_p2 = (deleted_zeros_32_fu_25545_p2 ^ 1'd1);

assign xor_ln895_71_fu_25591_p2 = (p_Result_103_reg_41396 ^ 1'd1);

assign xor_ln895_72_fu_25727_p2 = (deleted_zeros_33_fu_25692_p2 ^ 1'd1);

assign xor_ln895_73_fu_25739_p2 = (p_Result_106_reg_41427 ^ 1'd1);

assign xor_ln895_74_fu_25876_p2 = (deleted_zeros_34_fu_25841_p2 ^ 1'd1);

assign xor_ln895_75_fu_25888_p2 = (p_Result_109_reg_41456 ^ 1'd1);

assign xor_ln895_76_fu_26025_p2 = (deleted_zeros_35_fu_25990_p2 ^ 1'd1);

assign xor_ln895_77_fu_26037_p2 = (p_Result_112_reg_41485 ^ 1'd1);

assign xor_ln895_78_fu_22274_p2 = (deleted_zeros_36_fu_22236_p2 ^ 1'd1);

assign xor_ln895_79_fu_22286_p2 = (p_Result_115_fu_22148_p3 ^ 1'd1);

assign xor_ln895_7_fu_18825_p2 = (p_Result_9_reg_40400 ^ 1'd1);

assign xor_ln895_80_fu_26191_p2 = (deleted_zeros_37_fu_26156_p2 ^ 1'd1);

assign xor_ln895_81_fu_26203_p2 = (p_Result_118_reg_41529 ^ 1'd1);

assign xor_ln895_82_fu_26340_p2 = (deleted_zeros_38_fu_26305_p2 ^ 1'd1);

assign xor_ln895_83_fu_26352_p2 = (p_Result_121_reg_41558 ^ 1'd1);

assign xor_ln895_84_fu_26489_p2 = (deleted_zeros_39_fu_26454_p2 ^ 1'd1);

assign xor_ln895_85_fu_26501_p2 = (p_Result_124_reg_41587 ^ 1'd1);

assign xor_ln895_86_fu_26638_p2 = (deleted_zeros_40_fu_26603_p2 ^ 1'd1);

assign xor_ln895_87_fu_26650_p2 = (p_Result_127_reg_41616 ^ 1'd1);

assign xor_ln895_88_fu_26787_p2 = (deleted_zeros_41_fu_26752_p2 ^ 1'd1);

assign xor_ln895_89_fu_26799_p2 = (p_Result_130_reg_41645 ^ 1'd1);

assign xor_ln895_8_fu_18939_p2 = (deleted_zeros_4_fu_18904_p2 ^ 1'd1);

assign xor_ln895_90_fu_27010_p2 = (deleted_zeros_42_fu_26972_p2 ^ 1'd1);

assign xor_ln895_91_fu_27022_p2 = (p_Result_133_fu_26893_p3 ^ 1'd1);

assign xor_ln895_92_fu_30688_p2 = (deleted_zeros_43_fu_30653_p2 ^ 1'd1);

assign xor_ln895_93_fu_30699_p2 = (p_Result_136_reg_41771 ^ 1'd1);

assign xor_ln895_94_fu_30813_p2 = (deleted_zeros_44_fu_30778_p2 ^ 1'd1);

assign xor_ln895_95_fu_30824_p2 = (p_Result_139_reg_41802 ^ 1'd1);

assign xor_ln895_96_fu_30938_p2 = (deleted_zeros_45_fu_30903_p2 ^ 1'd1);

assign xor_ln895_97_fu_30949_p2 = (p_Result_142_reg_41833 ^ 1'd1);

assign xor_ln895_98_fu_31063_p2 = (deleted_zeros_46_fu_31028_p2 ^ 1'd1);

assign xor_ln895_99_fu_31074_p2 = (p_Result_145_reg_41864 ^ 1'd1);

assign xor_ln895_9_fu_18950_p2 = (p_Result_12_reg_40431 ^ 1'd1);

assign xor_ln895_fu_18547_p2 = (deleted_zeros_fu_18512_p2 ^ 1'd1);

assign xor_ln896_100_fu_31133_p2 = (p_Result_150_reg_41912 ^ 1'd1);

assign xor_ln896_101_fu_31210_p2 = (deleted_ones_50_fu_31178_p2 ^ 1'd1);

assign xor_ln896_102_fu_27474_p2 = (p_Result_153_fu_27466_p3 ^ 1'd1);

assign xor_ln896_103_fu_27568_p2 = (deleted_ones_51_fu_27532_p2 ^ 1'd1);

assign xor_ln896_104_fu_31275_p2 = (p_Result_156_reg_41958 ^ 1'd1);

assign xor_ln896_105_fu_31352_p2 = (deleted_ones_52_fu_31320_p2 ^ 1'd1);

assign xor_ln896_106_fu_27735_p2 = (p_Result_159_fu_27727_p3 ^ 1'd1);

assign xor_ln896_107_fu_27829_p2 = (deleted_ones_53_fu_27793_p2 ^ 1'd1);

assign xor_ln896_108_fu_31438_p2 = (p_Result_162_fu_31430_p3 ^ 1'd1);

assign xor_ln896_109_fu_31518_p2 = (deleted_ones_54_fu_31485_p2 ^ 1'd1);

assign xor_ln896_10_fu_19009_p2 = (p_Result_17_reg_40479 ^ 1'd1);

assign xor_ln896_110_fu_31587_p2 = (p_Result_165_fu_31579_p3 ^ 1'd1);

assign xor_ln896_111_fu_31667_p2 = (deleted_ones_55_fu_31634_p2 ^ 1'd1);

assign xor_ln896_112_fu_31736_p2 = (p_Result_168_fu_31728_p3 ^ 1'd1);

assign xor_ln896_113_fu_31816_p2 = (deleted_ones_56_fu_31783_p2 ^ 1'd1);

assign xor_ln896_114_fu_31885_p2 = (p_Result_171_fu_31877_p3 ^ 1'd1);

assign xor_ln896_115_fu_31965_p2 = (deleted_ones_57_fu_31932_p2 ^ 1'd1);

assign xor_ln896_116_fu_32034_p2 = (p_Result_174_fu_32026_p3 ^ 1'd1);

assign xor_ln896_117_fu_32114_p2 = (deleted_ones_58_fu_32081_p2 ^ 1'd1);

assign xor_ln896_118_fu_32183_p2 = (p_Result_177_fu_32175_p3 ^ 1'd1);

assign xor_ln896_119_fu_32263_p2 = (deleted_ones_59_fu_32230_p2 ^ 1'd1);

assign xor_ln896_11_fu_19086_p2 = (deleted_ones_5_fu_19054_p2 ^ 1'd1);

assign xor_ln896_120_fu_32332_p2 = (p_Result_180_fu_32324_p3 ^ 1'd1);

assign xor_ln896_121_fu_32412_p2 = (deleted_ones_60_fu_32379_p2 ^ 1'd1);

assign xor_ln896_122_fu_28257_p2 = (p_Result_183_fu_28249_p3 ^ 1'd1);

assign xor_ln896_123_fu_28351_p2 = (deleted_ones_61_fu_28315_p2 ^ 1'd1);

assign xor_ln896_124_fu_32498_p2 = (p_Result_186_fu_32490_p3 ^ 1'd1);

assign xor_ln896_125_fu_32578_p2 = (deleted_ones_62_fu_32545_p2 ^ 1'd1);

assign xor_ln896_126_fu_36163_p2 = (p_Result_189_reg_42403 ^ 1'd1);

assign xor_ln896_127_fu_36240_p2 = (deleted_ones_63_fu_36208_p2 ^ 1'd1);

assign xor_ln896_128_fu_36288_p2 = (p_Result_192_reg_42434 ^ 1'd1);

assign xor_ln896_129_fu_36365_p2 = (deleted_ones_64_fu_36333_p2 ^ 1'd1);

assign xor_ln896_12_fu_16881_p2 = (p_Result_20_fu_16873_p3 ^ 1'd1);

assign xor_ln896_130_fu_36413_p2 = (p_Result_195_reg_42465 ^ 1'd1);

assign xor_ln896_131_fu_36490_p2 = (deleted_ones_65_fu_36458_p2 ^ 1'd1);

assign xor_ln896_132_fu_36538_p2 = (p_Result_198_reg_42496 ^ 1'd1);

assign xor_ln896_133_fu_36615_p2 = (deleted_ones_66_fu_36583_p2 ^ 1'd1);

assign xor_ln896_134_fu_36663_p2 = (p_Result_201_reg_42527 ^ 1'd1);

assign xor_ln896_135_fu_36740_p2 = (deleted_ones_67_fu_36708_p2 ^ 1'd1);

assign xor_ln896_136_fu_33033_p2 = (p_Result_204_fu_33025_p3 ^ 1'd1);

assign xor_ln896_137_fu_33127_p2 = (deleted_ones_68_fu_33091_p2 ^ 1'd1);

assign xor_ln896_138_fu_36805_p2 = (p_Result_207_reg_42573 ^ 1'd1);

assign xor_ln896_139_fu_36882_p2 = (deleted_ones_69_fu_36850_p2 ^ 1'd1);

assign xor_ln896_13_fu_16975_p2 = (deleted_ones_6_fu_16939_p2 ^ 1'd1);

assign xor_ln896_140_fu_36930_p2 = (p_Result_210_reg_42604 ^ 1'd1);

assign xor_ln896_141_fu_37007_p2 = (deleted_ones_70_fu_36975_p2 ^ 1'd1);

assign xor_ln896_142_fu_37055_p2 = (p_Result_213_reg_42635 ^ 1'd1);

assign xor_ln896_143_fu_37132_p2 = (deleted_ones_71_fu_37100_p2 ^ 1'd1);

assign xor_ln896_144_fu_37201_p2 = (p_Result_216_fu_37193_p3 ^ 1'd1);

assign xor_ln896_145_fu_37281_p2 = (deleted_ones_72_fu_37248_p2 ^ 1'd1);

assign xor_ln896_146_fu_37350_p2 = (p_Result_219_fu_37342_p3 ^ 1'd1);

assign xor_ln896_147_fu_37430_p2 = (deleted_ones_73_fu_37397_p2 ^ 1'd1);

assign xor_ln896_148_fu_37499_p2 = (p_Result_222_fu_37491_p3 ^ 1'd1);

assign xor_ln896_149_fu_37579_p2 = (deleted_ones_74_fu_37546_p2 ^ 1'd1);

assign xor_ln896_14_fu_19148_p2 = (p_Result_23_reg_40525 ^ 1'd1);

assign xor_ln896_150_fu_37648_p2 = (p_Result_225_fu_37640_p3 ^ 1'd1);

assign xor_ln896_151_fu_37728_p2 = (deleted_ones_75_fu_37695_p2 ^ 1'd1);

assign xor_ln896_152_fu_33630_p2 = (p_Result_228_fu_33622_p3 ^ 1'd1);

assign xor_ln896_153_fu_33724_p2 = (deleted_ones_76_fu_33688_p2 ^ 1'd1);

assign xor_ln896_154_fu_37814_p2 = (p_Result_231_fu_37806_p3 ^ 1'd1);

assign xor_ln896_155_fu_37894_p2 = (deleted_ones_77_fu_37861_p2 ^ 1'd1);

assign xor_ln896_156_fu_37963_p2 = (p_Result_234_fu_37955_p3 ^ 1'd1);

assign xor_ln896_157_fu_38043_p2 = (deleted_ones_78_fu_38010_p2 ^ 1'd1);

assign xor_ln896_158_fu_38112_p2 = (p_Result_237_fu_38104_p3 ^ 1'd1);

assign xor_ln896_159_fu_38192_p2 = (deleted_ones_79_fu_38159_p2 ^ 1'd1);

assign xor_ln896_15_fu_19225_p2 = (deleted_ones_7_fu_19193_p2 ^ 1'd1);

assign xor_ln896_160_fu_38261_p2 = (p_Result_240_fu_38253_p3 ^ 1'd1);

assign xor_ln896_161_fu_38341_p2 = (deleted_ones_80_fu_38308_p2 ^ 1'd1);

assign xor_ln896_162_fu_22582_p2 = (p_Result_242_fu_22562_p3 ^ 1'd1);

assign xor_ln896_163_fu_22680_p2 = (p_Result_244_fu_22660_p3 ^ 1'd1);

assign xor_ln896_164_fu_22778_p2 = (p_Result_246_fu_22758_p3 ^ 1'd1);

assign xor_ln896_165_fu_22876_p2 = (p_Result_248_fu_22856_p3 ^ 1'd1);

assign xor_ln896_166_fu_22974_p2 = (p_Result_250_fu_22954_p3 ^ 1'd1);

assign xor_ln896_167_fu_23072_p2 = (p_Result_252_fu_23052_p3 ^ 1'd1);

assign xor_ln896_168_fu_23170_p2 = (p_Result_254_fu_23150_p3 ^ 1'd1);

assign xor_ln896_169_fu_23268_p2 = (p_Result_256_fu_23248_p3 ^ 1'd1);

assign xor_ln896_16_fu_19272_p2 = (p_Result_26_reg_40556 ^ 1'd1);

assign xor_ln896_170_fu_23366_p2 = (p_Result_258_fu_23346_p3 ^ 1'd1);

assign xor_ln896_171_fu_23468_p2 = (p_Result_260_fu_23448_p3 ^ 1'd1);

assign xor_ln896_172_fu_23570_p2 = (p_Result_262_fu_23550_p3 ^ 1'd1);

assign xor_ln896_173_fu_23672_p2 = (p_Result_264_fu_23652_p3 ^ 1'd1);

assign xor_ln896_174_fu_23774_p2 = (p_Result_266_fu_23754_p3 ^ 1'd1);

assign xor_ln896_175_fu_23876_p2 = (p_Result_268_fu_23856_p3 ^ 1'd1);

assign xor_ln896_176_fu_23978_p2 = (p_Result_270_fu_23958_p3 ^ 1'd1);

assign xor_ln896_177_fu_24080_p2 = (p_Result_272_fu_24060_p3 ^ 1'd1);

assign xor_ln896_178_fu_24182_p2 = (p_Result_274_fu_24162_p3 ^ 1'd1);

assign xor_ln896_179_fu_24284_p2 = (p_Result_276_fu_24264_p3 ^ 1'd1);

assign xor_ln896_17_fu_19349_p2 = (deleted_ones_8_fu_19317_p2 ^ 1'd1);

assign xor_ln896_180_fu_28469_p2 = (p_Result_278_fu_28449_p3 ^ 1'd1);

assign xor_ln896_181_fu_28569_p2 = (p_Result_280_fu_28549_p3 ^ 1'd1);

assign xor_ln896_182_fu_28633_p2 = (p_Result_282_reg_41729 ^ 1'd1);

assign xor_ln896_183_fu_28727_p2 = (p_Result_284_fu_28707_p3 ^ 1'd1);

assign xor_ln896_184_fu_28827_p2 = (p_Result_286_fu_28807_p3 ^ 1'd1);

assign xor_ln896_185_fu_28927_p2 = (p_Result_288_fu_28907_p3 ^ 1'd1);

assign xor_ln896_186_fu_28991_p2 = (p_Result_290_reg_41749 ^ 1'd1);

assign xor_ln896_187_fu_29085_p2 = (p_Result_292_fu_29065_p3 ^ 1'd1);

assign xor_ln896_188_fu_29185_p2 = (p_Result_294_fu_29165_p3 ^ 1'd1);

assign xor_ln896_189_fu_29287_p2 = (p_Result_296_fu_29267_p3 ^ 1'd1);

assign xor_ln896_18_fu_19418_p2 = (p_Result_29_fu_19410_p3 ^ 1'd1);

assign xor_ln896_190_fu_29389_p2 = (p_Result_298_fu_29369_p3 ^ 1'd1);

assign xor_ln896_191_fu_29491_p2 = (p_Result_300_fu_29471_p3 ^ 1'd1);

assign xor_ln896_192_fu_29593_p2 = (p_Result_302_fu_29573_p3 ^ 1'd1);

assign xor_ln896_193_fu_29695_p2 = (p_Result_304_fu_29675_p3 ^ 1'd1);

assign xor_ln896_194_fu_29797_p2 = (p_Result_306_fu_29777_p3 ^ 1'd1);

assign xor_ln896_195_fu_29899_p2 = (p_Result_308_fu_29879_p3 ^ 1'd1);

assign xor_ln896_196_fu_30001_p2 = (p_Result_310_fu_29981_p3 ^ 1'd1);

assign xor_ln896_197_fu_30103_p2 = (p_Result_312_fu_30083_p3 ^ 1'd1);

assign xor_ln896_198_fu_33932_p2 = (p_Result_314_reg_42247 ^ 1'd1);

assign xor_ln896_199_fu_33990_p2 = (p_Result_316_reg_42267 ^ 1'd1);

assign xor_ln896_19_fu_19498_p2 = (deleted_ones_9_fu_19465_p2 ^ 1'd1);

assign xor_ln896_1_fu_18569_p2 = (deleted_ones_fu_18537_p2 ^ 1'd1);

assign xor_ln896_200_fu_30277_p2 = (p_Result_318_fu_30257_p3 ^ 1'd1);

assign xor_ln896_201_fu_34048_p2 = (p_Result_320_reg_42293 ^ 1'd1);

assign xor_ln896_202_fu_34106_p2 = (p_Result_322_reg_42313 ^ 1'd1);

assign xor_ln896_203_fu_34164_p2 = (p_Result_324_reg_42333 ^ 1'd1);

assign xor_ln896_204_fu_30487_p2 = (p_Result_326_fu_30467_p3 ^ 1'd1);

assign xor_ln896_205_fu_34222_p2 = (p_Result_328_reg_42359 ^ 1'd1);

assign xor_ln896_206_fu_34280_p2 = (p_Result_330_reg_42379 ^ 1'd1);

assign xor_ln896_207_fu_34376_p2 = (p_Result_332_fu_34356_p3 ^ 1'd1);

assign xor_ln896_208_fu_34478_p2 = (p_Result_334_fu_34458_p3 ^ 1'd1);

assign xor_ln896_209_fu_34578_p2 = (p_Result_336_fu_34558_p3 ^ 1'd1);

assign xor_ln896_20_fu_17245_p2 = (p_Result_32_fu_17237_p3 ^ 1'd1);

assign xor_ln896_210_fu_34680_p2 = (p_Result_338_fu_34660_p3 ^ 1'd1);

assign xor_ln896_211_fu_34782_p2 = (p_Result_340_fu_34762_p3 ^ 1'd1);

assign xor_ln896_212_fu_34884_p2 = (p_Result_342_fu_34864_p3 ^ 1'd1);

assign xor_ln896_213_fu_34984_p2 = (p_Result_344_fu_34964_p3 ^ 1'd1);

assign xor_ln896_214_fu_35086_p2 = (p_Result_346_fu_35066_p3 ^ 1'd1);

assign xor_ln896_215_fu_35188_p2 = (p_Result_348_fu_35168_p3 ^ 1'd1);

assign xor_ln896_216_fu_35290_p2 = (p_Result_350_fu_35270_p3 ^ 1'd1);

assign xor_ln896_217_fu_35392_p2 = (p_Result_352_fu_35372_p3 ^ 1'd1);

assign xor_ln896_218_fu_35494_p2 = (p_Result_354_fu_35474_p3 ^ 1'd1);

assign xor_ln896_219_fu_35596_p2 = (p_Result_356_fu_35576_p3 ^ 1'd1);

assign xor_ln896_21_fu_17339_p2 = (deleted_ones_10_fu_17291_p2 ^ 1'd1);

assign xor_ln896_220_fu_35698_p2 = (p_Result_358_fu_35678_p3 ^ 1'd1);

assign xor_ln896_221_fu_35800_p2 = (p_Result_360_fu_35780_p3 ^ 1'd1);

assign xor_ln896_222_fu_35902_p2 = (p_Result_362_fu_35882_p3 ^ 1'd1);

assign xor_ln896_223_fu_36004_p2 = (p_Result_364_fu_35984_p3 ^ 1'd1);

assign xor_ln896_224_fu_36106_p2 = (p_Result_366_fu_36086_p3 ^ 1'd1);

assign xor_ln896_225_fu_38432_p2 = (p_Result_368_fu_38412_p3 ^ 1'd1);

assign xor_ln896_226_fu_38532_p2 = (p_Result_370_fu_38512_p3 ^ 1'd1);

assign xor_ln896_227_fu_38632_p2 = (p_Result_372_fu_38612_p3 ^ 1'd1);

assign xor_ln896_228_fu_38732_p2 = (p_Result_374_fu_38712_p3 ^ 1'd1);

assign xor_ln896_229_fu_38832_p2 = (p_Result_376_fu_38812_p3 ^ 1'd1);

assign xor_ln896_22_fu_17417_p2 = (p_Result_34_fu_17409_p3 ^ 1'd1);

assign xor_ln896_230_fu_38932_p2 = (p_Result_378_fu_38912_p3 ^ 1'd1);

assign xor_ln896_231_fu_39032_p2 = (p_Result_380_fu_39012_p3 ^ 1'd1);

assign xor_ln896_232_fu_39132_p2 = (p_Result_382_fu_39112_p3 ^ 1'd1);

assign xor_ln896_233_fu_39232_p2 = (p_Result_384_fu_39212_p3 ^ 1'd1);

assign xor_ln896_234_fu_39334_p2 = (p_Result_386_fu_39314_p3 ^ 1'd1);

assign xor_ln896_235_fu_39436_p2 = (p_Result_388_fu_39416_p3 ^ 1'd1);

assign xor_ln896_236_fu_39538_p2 = (p_Result_390_fu_39518_p3 ^ 1'd1);

assign xor_ln896_237_fu_39640_p2 = (p_Result_392_fu_39620_p3 ^ 1'd1);

assign xor_ln896_238_fu_39742_p2 = (p_Result_394_fu_39722_p3 ^ 1'd1);

assign xor_ln896_239_fu_39844_p2 = (p_Result_396_fu_39824_p3 ^ 1'd1);

assign xor_ln896_23_fu_17483_p2 = (deleted_ones_11_fu_17441_p2 ^ 1'd1);

assign xor_ln896_240_fu_39946_p2 = (p_Result_398_fu_39926_p3 ^ 1'd1);

assign xor_ln896_241_fu_40048_p2 = (p_Result_400_fu_40028_p3 ^ 1'd1);

assign xor_ln896_242_fu_40150_p2 = (p_Result_402_fu_40130_p3 ^ 1'd1);

assign xor_ln896_243_fu_18581_p2 = (or_ln896_fu_18575_p2 ^ and_ln891_fu_18542_p2);

assign xor_ln896_244_fu_18706_p2 = (or_ln896_1_fu_18700_p2 ^ and_ln891_1_fu_18667_p2);

assign xor_ln896_245_fu_16609_p2 = (or_ln896_2_fu_16603_p2 ^ and_ln891_2_fu_16567_p2);

assign xor_ln896_246_fu_18848_p2 = (or_ln896_3_fu_18842_p2 ^ and_ln891_3_fu_18809_p2);

assign xor_ln896_247_fu_18973_p2 = (or_ln896_4_fu_18967_p2 ^ and_ln891_4_fu_18934_p2);

assign xor_ln896_248_fu_19098_p2 = (or_ln896_5_fu_19092_p2 ^ and_ln891_5_fu_19059_p2);

assign xor_ln896_249_fu_16987_p2 = (or_ln896_6_fu_16981_p2 ^ and_ln891_6_fu_16945_p2);

assign xor_ln896_24_fu_19601_p2 = (p_Result_37_fu_19593_p3 ^ 1'd1);

assign xor_ln896_250_fu_19237_p2 = (or_ln896_7_fu_19231_p2 ^ and_ln891_7_fu_19198_p2);

assign xor_ln896_251_fu_19361_p2 = (or_ln896_8_fu_19355_p2 ^ and_ln891_8_fu_19322_p2);

assign xor_ln896_252_fu_19510_p2 = (or_ln896_9_fu_19504_p2 ^ and_ln891_9_fu_19470_p2);

assign xor_ln896_253_fu_17351_p2 = (or_ln896_10_fu_17345_p2 ^ and_ln891_10_fu_17303_p2);

assign xor_ln896_254_fu_17495_p2 = (or_ln896_11_fu_17489_p2 ^ and_ln891_11_fu_17453_p2);

assign xor_ln896_255_fu_19693_p2 = (or_ln896_12_fu_19687_p2 ^ and_ln891_12_fu_19653_p2);

assign xor_ln896_256_fu_19842_p2 = (or_ln896_13_fu_19836_p2 ^ and_ln891_13_fu_19802_p2);

assign xor_ln896_257_fu_17723_p2 = (or_ln896_14_fu_17717_p2 ^ and_ln891_14_fu_17681_p2);

assign xor_ln896_258_fu_19984_p2 = (or_ln896_15_fu_19978_p2 ^ and_ln891_15_fu_19945_p2);

assign xor_ln896_259_fu_20133_p2 = (or_ln896_16_fu_20127_p2 ^ and_ln891_16_fu_20093_p2);

assign xor_ln896_25_fu_19681_p2 = (deleted_ones_12_fu_19648_p2 ^ 1'd1);

assign xor_ln896_260_fu_20282_p2 = (or_ln896_17_fu_20276_p2 ^ and_ln891_17_fu_20242_p2);

assign xor_ln896_261_fu_20427_p2 = (or_ln896_18_fu_20421_p2 ^ and_ln891_18_fu_20387_p2);

assign xor_ln896_262_fu_20556_p2 = (or_ln896_19_fu_20550_p2 ^ and_ln891_19_fu_20516_p2);

assign xor_ln896_263_fu_20689_p2 = (or_ln896_20_fu_20683_p2 ^ and_ln891_20_fu_20649_p2);

assign xor_ln896_264_fu_20834_p2 = (or_ln896_21_fu_20828_p2 ^ and_ln891_21_fu_20794_p2);

assign xor_ln896_265_fu_20963_p2 = (or_ln896_22_fu_20957_p2 ^ and_ln891_22_fu_20923_p2);

assign xor_ln896_266_fu_21092_p2 = (or_ln896_23_fu_21086_p2 ^ and_ln891_23_fu_21052_p2);

assign xor_ln896_267_fu_18361_p2 = (or_ln896_24_fu_18355_p2 ^ and_ln891_24_fu_18319_p2);

assign xor_ln896_268_fu_21238_p2 = (or_ln896_25_fu_21232_p2 ^ and_ln891_25_fu_21198_p2);

assign xor_ln896_269_fu_21367_p2 = (or_ln896_26_fu_21361_p2 ^ and_ln891_26_fu_21327_p2);

assign xor_ln896_26_fu_19750_p2 = (p_Result_40_fu_19742_p3 ^ 1'd1);

assign xor_ln896_270_fu_24618_p2 = (or_ln896_27_fu_24612_p2 ^ and_ln891_27_fu_24579_p2);

assign xor_ln896_271_fu_24742_p2 = (or_ln896_28_fu_24736_p2 ^ and_ln891_28_fu_24703_p2);

assign xor_ln896_272_fu_24867_p2 = (or_ln896_29_fu_24861_p2 ^ and_ln891_29_fu_24828_p2);

assign xor_ln896_273_fu_24992_p2 = (or_ln896_30_fu_24986_p2 ^ and_ln891_30_fu_24953_p2);

assign xor_ln896_274_fu_25117_p2 = (or_ln896_31_fu_25111_p2 ^ and_ln891_31_fu_25078_p2);

assign xor_ln896_275_fu_25242_p2 = (or_ln896_32_fu_25236_p2 ^ and_ln891_32_fu_25203_p2);

assign xor_ln896_276_fu_25367_p2 = (or_ln896_33_fu_25361_p2 ^ and_ln891_33_fu_25328_p2);

assign xor_ln896_277_fu_25492_p2 = (or_ln896_34_fu_25486_p2 ^ and_ln891_34_fu_25453_p2);

assign xor_ln896_278_fu_25614_p2 = (or_ln896_35_fu_25608_p2 ^ and_ln891_35_fu_25575_p2);

assign xor_ln896_279_fu_25762_p2 = (or_ln896_36_fu_25756_p2 ^ and_ln891_36_fu_25722_p2);

assign xor_ln896_27_fu_19830_p2 = (deleted_ones_13_fu_19797_p2 ^ 1'd1);

assign xor_ln896_280_fu_25911_p2 = (or_ln896_37_fu_25905_p2 ^ and_ln891_37_fu_25871_p2);

assign xor_ln896_281_fu_26060_p2 = (or_ln896_38_fu_26054_p2 ^ and_ln891_38_fu_26020_p2);

assign xor_ln896_282_fu_22310_p2 = (or_ln896_39_fu_22304_p2 ^ and_ln891_39_fu_22268_p2);

assign xor_ln896_283_fu_26226_p2 = (or_ln896_40_fu_26220_p2 ^ and_ln891_40_fu_26186_p2);

assign xor_ln896_284_fu_26375_p2 = (or_ln896_41_fu_26369_p2 ^ and_ln891_41_fu_26335_p2);

assign xor_ln896_285_fu_26524_p2 = (or_ln896_42_fu_26518_p2 ^ and_ln891_42_fu_26484_p2);

assign xor_ln896_286_fu_26673_p2 = (or_ln896_43_fu_26667_p2 ^ and_ln891_43_fu_26633_p2);

assign xor_ln896_287_fu_26822_p2 = (or_ln896_44_fu_26816_p2 ^ and_ln891_44_fu_26782_p2);

assign xor_ln896_288_fu_27046_p2 = (or_ln896_45_fu_27040_p2 ^ and_ln891_45_fu_27004_p2);

assign xor_ln896_289_fu_30722_p2 = (or_ln896_46_fu_30716_p2 ^ and_ln891_46_fu_30683_p2);

assign xor_ln896_28_fu_17645_p2 = (p_Result_42_fu_17637_p3 ^ 1'd1);

assign xor_ln896_290_fu_30847_p2 = (or_ln896_47_fu_30841_p2 ^ and_ln891_47_fu_30808_p2);

assign xor_ln896_291_fu_30972_p2 = (or_ln896_48_fu_30966_p2 ^ and_ln891_48_fu_30933_p2);

assign xor_ln896_292_fu_31097_p2 = (or_ln896_49_fu_31091_p2 ^ and_ln891_49_fu_31058_p2);

assign xor_ln896_293_fu_31222_p2 = (or_ln896_50_fu_31216_p2 ^ and_ln891_50_fu_31183_p2);

assign xor_ln896_294_fu_27580_p2 = (or_ln896_51_fu_27574_p2 ^ and_ln891_51_fu_27538_p2);

assign xor_ln896_295_fu_31364_p2 = (or_ln896_52_fu_31358_p2 ^ and_ln891_52_fu_31325_p2);

assign xor_ln896_296_fu_27841_p2 = (or_ln896_53_fu_27835_p2 ^ and_ln891_53_fu_27799_p2);

assign xor_ln896_297_fu_31530_p2 = (or_ln896_54_fu_31524_p2 ^ and_ln891_54_fu_31490_p2);

assign xor_ln896_298_fu_31679_p2 = (or_ln896_55_fu_31673_p2 ^ and_ln891_55_fu_31639_p2);

assign xor_ln896_299_fu_31828_p2 = (or_ln896_56_fu_31822_p2 ^ and_ln891_56_fu_31788_p2);

assign xor_ln896_29_fu_17711_p2 = (deleted_ones_14_fu_17669_p2 ^ 1'd1);

assign xor_ln896_2_fu_18617_p2 = (p_Result_5_reg_40371 ^ 1'd1);

assign xor_ln896_300_fu_31977_p2 = (or_ln896_57_fu_31971_p2 ^ and_ln891_57_fu_31937_p2);

assign xor_ln896_301_fu_32126_p2 = (or_ln896_58_fu_32120_p2 ^ and_ln891_58_fu_32086_p2);

assign xor_ln896_302_fu_32275_p2 = (or_ln896_59_fu_32269_p2 ^ and_ln891_59_fu_32235_p2);

assign xor_ln896_303_fu_32424_p2 = (or_ln896_60_fu_32418_p2 ^ and_ln891_60_fu_32384_p2);

assign xor_ln896_304_fu_28363_p2 = (or_ln896_61_fu_28357_p2 ^ and_ln891_61_fu_28321_p2);

assign xor_ln896_305_fu_32590_p2 = (or_ln896_62_fu_32584_p2 ^ and_ln891_62_fu_32550_p2);

assign xor_ln896_306_fu_36252_p2 = (or_ln896_63_fu_36246_p2 ^ and_ln891_63_fu_36213_p2);

assign xor_ln896_307_fu_36377_p2 = (or_ln896_64_fu_36371_p2 ^ and_ln891_64_fu_36338_p2);

assign xor_ln896_308_fu_36502_p2 = (or_ln896_65_fu_36496_p2 ^ and_ln891_65_fu_36463_p2);

assign xor_ln896_309_fu_36627_p2 = (or_ln896_66_fu_36621_p2 ^ and_ln891_66_fu_36588_p2);

assign xor_ln896_30_fu_19895_p2 = (p_Result_45_reg_40719 ^ 1'd1);

assign xor_ln896_310_fu_36752_p2 = (or_ln896_67_fu_36746_p2 ^ and_ln891_67_fu_36713_p2);

assign xor_ln896_311_fu_33139_p2 = (or_ln896_68_fu_33133_p2 ^ and_ln891_68_fu_33097_p2);

assign xor_ln896_312_fu_36894_p2 = (or_ln896_69_fu_36888_p2 ^ and_ln891_69_fu_36855_p2);

assign xor_ln896_313_fu_37019_p2 = (or_ln896_70_fu_37013_p2 ^ and_ln891_70_fu_36980_p2);

assign xor_ln896_314_fu_37144_p2 = (or_ln896_71_fu_37138_p2 ^ and_ln891_71_fu_37105_p2);

assign xor_ln896_315_fu_37293_p2 = (or_ln896_72_fu_37287_p2 ^ and_ln891_72_fu_37253_p2);

assign xor_ln896_316_fu_37442_p2 = (or_ln896_73_fu_37436_p2 ^ and_ln891_73_fu_37402_p2);

assign xor_ln896_317_fu_37591_p2 = (or_ln896_74_fu_37585_p2 ^ and_ln891_74_fu_37551_p2);

assign xor_ln896_318_fu_37740_p2 = (or_ln896_75_fu_37734_p2 ^ and_ln891_75_fu_37700_p2);

assign xor_ln896_319_fu_33736_p2 = (or_ln896_76_fu_33730_p2 ^ and_ln891_76_fu_33694_p2);

assign xor_ln896_31_fu_19972_p2 = (deleted_ones_15_fu_19940_p2 ^ 1'd1);

assign xor_ln896_320_fu_37906_p2 = (or_ln896_77_fu_37900_p2 ^ and_ln891_77_fu_37866_p2);

assign xor_ln896_321_fu_38055_p2 = (or_ln896_78_fu_38049_p2 ^ and_ln891_78_fu_38015_p2);

assign xor_ln896_322_fu_38204_p2 = (or_ln896_79_fu_38198_p2 ^ and_ln891_79_fu_38164_p2);

assign xor_ln896_323_fu_38353_p2 = (or_ln896_80_fu_38347_p2 ^ and_ln891_80_fu_38313_p2);

assign xor_ln896_32_fu_20041_p2 = (p_Result_48_fu_20033_p3 ^ 1'd1);

assign xor_ln896_33_fu_20121_p2 = (deleted_ones_16_fu_20088_p2 ^ 1'd1);

assign xor_ln896_34_fu_20190_p2 = (p_Result_51_fu_20182_p3 ^ 1'd1);

assign xor_ln896_35_fu_20270_p2 = (deleted_ones_17_fu_20237_p2 ^ 1'd1);

assign xor_ln896_36_fu_20335_p2 = (p_Result_54_fu_20327_p3 ^ 1'd1);

assign xor_ln896_37_fu_20415_p2 = (deleted_ones_18_fu_20382_p2 ^ 1'd1);

assign xor_ln896_38_fu_20464_p2 = (p_Result_57_fu_20456_p3 ^ 1'd1);

assign xor_ln896_39_fu_20544_p2 = (deleted_ones_19_fu_20511_p2 ^ 1'd1);

assign xor_ln896_3_fu_18694_p2 = (deleted_ones_1_fu_18662_p2 ^ 1'd1);

assign xor_ln896_40_fu_20597_p2 = (p_Result_60_fu_20589_p3 ^ 1'd1);

assign xor_ln896_41_fu_20677_p2 = (deleted_ones_20_fu_20644_p2 ^ 1'd1);

assign xor_ln896_42_fu_20742_p2 = (p_Result_63_fu_20734_p3 ^ 1'd1);

assign xor_ln896_43_fu_20822_p2 = (deleted_ones_21_fu_20789_p2 ^ 1'd1);

assign xor_ln896_44_fu_20871_p2 = (p_Result_66_fu_20863_p3 ^ 1'd1);

assign xor_ln896_45_fu_20951_p2 = (deleted_ones_22_fu_20918_p2 ^ 1'd1);

assign xor_ln896_46_fu_21000_p2 = (p_Result_69_fu_20992_p3 ^ 1'd1);

assign xor_ln896_47_fu_21080_p2 = (deleted_ones_23_fu_21047_p2 ^ 1'd1);

assign xor_ln896_48_fu_18255_p2 = (p_Result_72_fu_18247_p3 ^ 1'd1);

assign xor_ln896_49_fu_18349_p2 = (deleted_ones_24_fu_18313_p2 ^ 1'd1);

assign xor_ln896_4_fu_16503_p2 = (p_Result_8_fu_16495_p3 ^ 1'd1);

assign xor_ln896_50_fu_21146_p2 = (p_Result_75_fu_21138_p3 ^ 1'd1);

assign xor_ln896_51_fu_21226_p2 = (deleted_ones_25_fu_21193_p2 ^ 1'd1);

assign xor_ln896_52_fu_21275_p2 = (p_Result_78_fu_21267_p3 ^ 1'd1);

assign xor_ln896_53_fu_21355_p2 = (deleted_ones_26_fu_21322_p2 ^ 1'd1);

assign xor_ln896_54_fu_24529_p2 = (p_Result_81_reg_41165 ^ 1'd1);

assign xor_ln896_55_fu_24606_p2 = (deleted_ones_27_fu_24574_p2 ^ 1'd1);

assign xor_ln896_56_fu_24653_p2 = (p_Result_84_reg_41196 ^ 1'd1);

assign xor_ln896_57_fu_24730_p2 = (deleted_ones_28_fu_24698_p2 ^ 1'd1);

assign xor_ln896_58_fu_24778_p2 = (p_Result_87_reg_41227 ^ 1'd1);

assign xor_ln896_59_fu_24855_p2 = (deleted_ones_29_fu_24823_p2 ^ 1'd1);

assign xor_ln896_5_fu_16597_p2 = (deleted_ones_2_fu_16561_p2 ^ 1'd1);

assign xor_ln896_60_fu_24903_p2 = (p_Result_90_reg_41258 ^ 1'd1);

assign xor_ln896_61_fu_24980_p2 = (deleted_ones_30_fu_24948_p2 ^ 1'd1);

assign xor_ln896_62_fu_25028_p2 = (p_Result_93_reg_41289 ^ 1'd1);

assign xor_ln896_63_fu_25105_p2 = (deleted_ones_31_fu_25073_p2 ^ 1'd1);

assign xor_ln896_64_fu_25153_p2 = (p_Result_96_reg_41320 ^ 1'd1);

assign xor_ln896_65_fu_25230_p2 = (deleted_ones_32_fu_25198_p2 ^ 1'd1);

assign xor_ln896_66_fu_25278_p2 = (p_Result_99_reg_41351 ^ 1'd1);

assign xor_ln896_67_fu_25355_p2 = (deleted_ones_33_fu_25323_p2 ^ 1'd1);

assign xor_ln896_68_fu_25403_p2 = (p_Result_102_reg_41382 ^ 1'd1);

assign xor_ln896_69_fu_25480_p2 = (deleted_ones_34_fu_25448_p2 ^ 1'd1);

assign xor_ln896_6_fu_18759_p2 = (p_Result_11_reg_40417 ^ 1'd1);

assign xor_ln896_70_fu_25525_p2 = (p_Result_105_reg_41413 ^ 1'd1);

assign xor_ln896_71_fu_25602_p2 = (deleted_ones_35_fu_25570_p2 ^ 1'd1);

assign xor_ln896_72_fu_25670_p2 = (p_Result_108_fu_25662_p3 ^ 1'd1);

assign xor_ln896_73_fu_25750_p2 = (deleted_ones_36_fu_25717_p2 ^ 1'd1);

assign xor_ln896_74_fu_25819_p2 = (p_Result_111_fu_25811_p3 ^ 1'd1);

assign xor_ln896_75_fu_25899_p2 = (deleted_ones_37_fu_25866_p2 ^ 1'd1);

assign xor_ln896_76_fu_25968_p2 = (p_Result_114_fu_25960_p3 ^ 1'd1);

assign xor_ln896_77_fu_26048_p2 = (deleted_ones_38_fu_26015_p2 ^ 1'd1);

assign xor_ln896_78_fu_22204_p2 = (p_Result_117_fu_22196_p3 ^ 1'd1);

assign xor_ln896_79_fu_22298_p2 = (deleted_ones_39_fu_22262_p2 ^ 1'd1);

assign xor_ln896_7_fu_18836_p2 = (deleted_ones_3_fu_18804_p2 ^ 1'd1);

assign xor_ln896_80_fu_26134_p2 = (p_Result_120_fu_26126_p3 ^ 1'd1);

assign xor_ln896_81_fu_26214_p2 = (deleted_ones_40_fu_26181_p2 ^ 1'd1);

assign xor_ln896_82_fu_26283_p2 = (p_Result_123_fu_26275_p3 ^ 1'd1);

assign xor_ln896_83_fu_26363_p2 = (deleted_ones_41_fu_26330_p2 ^ 1'd1);

assign xor_ln896_84_fu_26432_p2 = (p_Result_126_fu_26424_p3 ^ 1'd1);

assign xor_ln896_85_fu_26512_p2 = (deleted_ones_42_fu_26479_p2 ^ 1'd1);

assign xor_ln896_86_fu_26581_p2 = (p_Result_129_fu_26573_p3 ^ 1'd1);

assign xor_ln896_87_fu_26661_p2 = (deleted_ones_43_fu_26628_p2 ^ 1'd1);

assign xor_ln896_88_fu_26730_p2 = (p_Result_132_fu_26722_p3 ^ 1'd1);

assign xor_ln896_89_fu_26810_p2 = (deleted_ones_44_fu_26777_p2 ^ 1'd1);

assign xor_ln896_8_fu_18884_p2 = (p_Result_14_reg_40448 ^ 1'd1);

assign xor_ln896_90_fu_26940_p2 = (p_Result_135_fu_26932_p3 ^ 1'd1);

assign xor_ln896_91_fu_27034_p2 = (deleted_ones_45_fu_26998_p2 ^ 1'd1);

assign xor_ln896_92_fu_30633_p2 = (p_Result_138_reg_41788 ^ 1'd1);

assign xor_ln896_93_fu_30710_p2 = (deleted_ones_46_fu_30678_p2 ^ 1'd1);

assign xor_ln896_94_fu_30758_p2 = (p_Result_141_reg_41819 ^ 1'd1);

assign xor_ln896_95_fu_30835_p2 = (deleted_ones_47_fu_30803_p2 ^ 1'd1);

assign xor_ln896_96_fu_30883_p2 = (p_Result_144_reg_41850 ^ 1'd1);

assign xor_ln896_97_fu_30960_p2 = (deleted_ones_48_fu_30928_p2 ^ 1'd1);

assign xor_ln896_98_fu_31008_p2 = (p_Result_147_reg_41881 ^ 1'd1);

assign xor_ln896_99_fu_31085_p2 = (deleted_ones_49_fu_31053_p2 ^ 1'd1);

assign xor_ln896_9_fu_18961_p2 = (deleted_ones_4_fu_18929_p2 ^ 1'd1);

assign xor_ln896_fu_18492_p2 = (p_Result_2_reg_40340 ^ 1'd1);

assign zext_ln377_10_fu_17227_p1 = tmp_60_fu_17219_p3;

assign zext_ln377_11_fu_17399_p1 = tmp_65_fu_17391_p3;

assign zext_ln377_12_fu_19580_p1 = tmp_69_reg_40646;

assign zext_ln377_13_fu_19729_p1 = tmp_75_reg_40675;

assign zext_ln377_14_fu_17627_p1 = tmp_80_fu_17619_p3;

assign zext_ln377_15_fu_17779_p1 = tmp_84_fu_17771_p3;

assign zext_ln377_16_fu_20020_p1 = tmp_90_reg_40750;

assign zext_ln377_17_fu_20169_p1 = tmp_96_reg_40779;

assign zext_ln377_18_fu_20318_p1 = tmp_102_reg_40808;

assign zext_ln377_19_fu_20447_p1 = tmp_108_reg_40837;

assign zext_ln377_1_fu_16385_p1 = tmp_6_fu_16377_p3;

assign zext_ln377_20_fu_20576_p1 = tmp_114_reg_40866;

assign zext_ln377_21_fu_20725_p1 = tmp_120_reg_40895;

assign zext_ln377_22_fu_20854_p1 = tmp_126_reg_40924;

assign zext_ln377_23_fu_20983_p1 = tmp_132_reg_40953;

assign zext_ln377_24_fu_18237_p1 = tmp_138_fu_18229_p3;

assign zext_ln377_25_fu_21129_p1 = tmp_144_reg_40997;

assign zext_ln377_26_fu_21258_p1 = tmp_150_reg_41026;

assign zext_ln377_27_fu_21442_p1 = tmp_156_fu_21434_p3;

assign zext_ln377_28_fu_21506_p1 = tmp_162_fu_21498_p3;

assign zext_ln377_29_fu_21570_p1 = tmp_168_fu_21562_p3;

assign zext_ln377_2_fu_16485_p1 = tmp_12_fu_16477_p3;

assign zext_ln377_30_fu_21634_p1 = tmp_174_fu_21626_p3;

assign zext_ln377_31_fu_21698_p1 = tmp_180_fu_21690_p3;

assign zext_ln377_32_fu_21762_p1 = tmp_186_fu_21754_p3;

assign zext_ln377_33_fu_21826_p1 = tmp_192_fu_21818_p3;

assign zext_ln377_34_fu_21890_p1 = tmp_198_fu_21882_p3;

assign zext_ln377_35_fu_21950_p1 = tmp_204_fu_21942_p3;

assign zext_ln377_36_fu_25649_p1 = tmp_210_reg_41444;

assign zext_ln377_37_fu_25798_p1 = tmp_216_reg_41473;

assign zext_ln377_38_fu_25947_p1 = tmp_222_reg_41502;

assign zext_ln377_39_fu_22186_p1 = tmp_228_fu_22178_p3;

assign zext_ln377_3_fu_16665_p1 = tmp_18_fu_16657_p3;

assign zext_ln377_40_fu_26113_p1 = tmp_234_reg_41546;

assign zext_ln377_41_fu_26262_p1 = tmp_240_reg_41575;

assign zext_ln377_42_fu_26411_p1 = tmp_246_reg_41604;

assign zext_ln377_43_fu_26560_p1 = tmp_252_reg_41633;

assign zext_ln377_44_fu_26709_p1 = tmp_258_reg_41662;

assign zext_ln377_45_fu_26923_p1 = tmp_264_reg_41038_pp0_iter1_reg;

assign zext_ln377_46_fu_27102_p1 = tmp_270_fu_27094_p3;

assign zext_ln377_47_fu_27166_p1 = tmp_276_fu_27158_p3;

assign zext_ln377_48_fu_27230_p1 = tmp_282_fu_27222_p3;

assign zext_ln377_49_fu_27294_p1 = tmp_288_fu_27286_p3;

assign zext_ln377_4_fu_16729_p1 = tmp_24_fu_16721_p3;

assign zext_ln377_50_fu_27358_p1 = tmp_294_fu_27350_p3;

assign zext_ln377_51_fu_27456_p1 = tmp_300_fu_27448_p3;

assign zext_ln377_52_fu_27636_p1 = tmp_306_fu_27628_p3;

assign zext_ln377_53_fu_27717_p1 = tmp_312_fu_27709_p3;

assign zext_ln377_54_fu_31417_p1 = tmp_318_reg_42004;

assign zext_ln377_55_fu_31566_p1 = tmp_324_reg_42033;

assign zext_ln377_56_fu_31715_p1 = tmp_330_reg_42062;

assign zext_ln377_57_fu_31864_p1 = tmp_336_reg_42091;

assign zext_ln377_58_fu_32013_p1 = tmp_342_reg_42120;

assign zext_ln377_59_fu_32162_p1 = tmp_348_reg_42149;

assign zext_ln377_5_fu_16793_p1 = tmp_30_fu_16785_p3;

assign zext_ln377_60_fu_32311_p1 = tmp_354_reg_42178;

assign zext_ln377_61_fu_28239_p1 = tmp_360_fu_28231_p3;

assign zext_ln377_62_fu_32477_p1 = tmp_366_reg_42222;

assign zext_ln377_63_fu_32678_p1 = tmp_372_fu_32670_p3;

assign zext_ln377_64_fu_32742_p1 = tmp_378_fu_32734_p3;

assign zext_ln377_65_fu_32806_p1 = tmp_384_fu_32798_p3;

assign zext_ln377_66_fu_32870_p1 = tmp_390_fu_32862_p3;

assign zext_ln377_67_fu_32934_p1 = tmp_396_fu_32926_p3;

assign zext_ln377_68_fu_33015_p1 = tmp_402_fu_33007_p3;

assign zext_ln377_69_fu_33195_p1 = tmp_408_fu_33187_p3;

assign zext_ln377_6_fu_16863_p1 = tmp_36_fu_16855_p3;

assign zext_ln377_70_fu_33259_p1 = tmp_414_fu_33251_p3;

assign zext_ln377_71_fu_33323_p1 = tmp_420_fu_33315_p3;

assign zext_ln377_72_fu_37180_p1 = tmp_426_reg_42666;

assign zext_ln377_73_fu_37329_p1 = tmp_432_reg_42695;

assign zext_ln377_74_fu_37478_p1 = tmp_438_reg_42724;

assign zext_ln377_75_fu_37627_p1 = tmp_444_reg_42753;

assign zext_ln377_76_fu_33612_p1 = tmp_450_fu_33604_p3;

assign zext_ln377_77_fu_37793_p1 = tmp_456_reg_42797;

assign zext_ln377_78_fu_37942_p1 = tmp_462_reg_42826;

assign zext_ln377_79_fu_38091_p1 = tmp_468_reg_42855;

assign zext_ln377_7_fu_17039_p1 = tmp_42_fu_17031_p3;

assign zext_ln377_80_fu_38240_p1 = tmp_474_reg_42884;

assign zext_ln377_8_fu_17103_p1 = tmp_48_fu_17095_p3;

assign zext_ln377_9_fu_19397_p1 = tmp_54_reg_40587;

assign zext_ln377_fu_16321_p1 = tmp_fu_16313_p3;

endmodule //motorB_dense_latency_ap_fixed_32_8_0_0_0_ap_fixed_32_8_0_0_0_config8_s
