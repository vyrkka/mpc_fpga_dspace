module mpc_qp_admm (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        p_read2,
        h_address0,
        h_ce0,
        h_q0,
        h_address1,
        h_ce1,
        h_q1,
        xk_admm_V_0,
        xk_admm_V_0_ap_vld
);

parameter    ap_ST_fsm_state1 = 85'd1;
parameter    ap_ST_fsm_state2 = 85'd2;
parameter    ap_ST_fsm_state3 = 85'd4;
parameter    ap_ST_fsm_state4 = 85'd8;
parameter    ap_ST_fsm_state5 = 85'd16;
parameter    ap_ST_fsm_state6 = 85'd32;
parameter    ap_ST_fsm_state7 = 85'd64;
parameter    ap_ST_fsm_state8 = 85'd128;
parameter    ap_ST_fsm_state9 = 85'd256;
parameter    ap_ST_fsm_state10 = 85'd512;
parameter    ap_ST_fsm_state11 = 85'd1024;
parameter    ap_ST_fsm_state12 = 85'd2048;
parameter    ap_ST_fsm_state13 = 85'd4096;
parameter    ap_ST_fsm_state14 = 85'd8192;
parameter    ap_ST_fsm_state15 = 85'd16384;
parameter    ap_ST_fsm_state16 = 85'd32768;
parameter    ap_ST_fsm_state17 = 85'd65536;
parameter    ap_ST_fsm_state18 = 85'd131072;
parameter    ap_ST_fsm_state19 = 85'd262144;
parameter    ap_ST_fsm_state20 = 85'd524288;
parameter    ap_ST_fsm_state21 = 85'd1048576;
parameter    ap_ST_fsm_state22 = 85'd2097152;
parameter    ap_ST_fsm_state23 = 85'd4194304;
parameter    ap_ST_fsm_state24 = 85'd8388608;
parameter    ap_ST_fsm_state25 = 85'd16777216;
parameter    ap_ST_fsm_state26 = 85'd33554432;
parameter    ap_ST_fsm_state27 = 85'd67108864;
parameter    ap_ST_fsm_state28 = 85'd134217728;
parameter    ap_ST_fsm_state29 = 85'd268435456;
parameter    ap_ST_fsm_state30 = 85'd536870912;
parameter    ap_ST_fsm_state31 = 85'd1073741824;
parameter    ap_ST_fsm_state32 = 85'd2147483648;
parameter    ap_ST_fsm_state33 = 85'd4294967296;
parameter    ap_ST_fsm_state34 = 85'd8589934592;
parameter    ap_ST_fsm_state35 = 85'd17179869184;
parameter    ap_ST_fsm_state36 = 85'd34359738368;
parameter    ap_ST_fsm_state37 = 85'd68719476736;
parameter    ap_ST_fsm_state38 = 85'd137438953472;
parameter    ap_ST_fsm_state39 = 85'd274877906944;
parameter    ap_ST_fsm_state40 = 85'd549755813888;
parameter    ap_ST_fsm_state41 = 85'd1099511627776;
parameter    ap_ST_fsm_state42 = 85'd2199023255552;
parameter    ap_ST_fsm_state43 = 85'd4398046511104;
parameter    ap_ST_fsm_state44 = 85'd8796093022208;
parameter    ap_ST_fsm_state45 = 85'd17592186044416;
parameter    ap_ST_fsm_state46 = 85'd35184372088832;
parameter    ap_ST_fsm_state47 = 85'd70368744177664;
parameter    ap_ST_fsm_state48 = 85'd140737488355328;
parameter    ap_ST_fsm_state49 = 85'd281474976710656;
parameter    ap_ST_fsm_state50 = 85'd562949953421312;
parameter    ap_ST_fsm_state51 = 85'd1125899906842624;
parameter    ap_ST_fsm_state52 = 85'd2251799813685248;
parameter    ap_ST_fsm_state53 = 85'd4503599627370496;
parameter    ap_ST_fsm_state54 = 85'd9007199254740992;
parameter    ap_ST_fsm_state55 = 85'd18014398509481984;
parameter    ap_ST_fsm_state56 = 85'd36028797018963968;
parameter    ap_ST_fsm_state57 = 85'd72057594037927936;
parameter    ap_ST_fsm_state58 = 85'd144115188075855872;
parameter    ap_ST_fsm_state59 = 85'd288230376151711744;
parameter    ap_ST_fsm_state60 = 85'd576460752303423488;
parameter    ap_ST_fsm_state61 = 85'd1152921504606846976;
parameter    ap_ST_fsm_state62 = 85'd2305843009213693952;
parameter    ap_ST_fsm_state63 = 85'd4611686018427387904;
parameter    ap_ST_fsm_state64 = 85'd9223372036854775808;
parameter    ap_ST_fsm_state65 = 85'd18446744073709551616;
parameter    ap_ST_fsm_state66 = 85'd36893488147419103232;
parameter    ap_ST_fsm_state67 = 85'd73786976294838206464;
parameter    ap_ST_fsm_state68 = 85'd147573952589676412928;
parameter    ap_ST_fsm_state69 = 85'd295147905179352825856;
parameter    ap_ST_fsm_state70 = 85'd590295810358705651712;
parameter    ap_ST_fsm_state71 = 85'd1180591620717411303424;
parameter    ap_ST_fsm_state72 = 85'd2361183241434822606848;
parameter    ap_ST_fsm_state73 = 85'd4722366482869645213696;
parameter    ap_ST_fsm_state74 = 85'd9444732965739290427392;
parameter    ap_ST_fsm_state75 = 85'd18889465931478580854784;
parameter    ap_ST_fsm_state76 = 85'd37778931862957161709568;
parameter    ap_ST_fsm_state77 = 85'd75557863725914323419136;
parameter    ap_ST_fsm_state78 = 85'd151115727451828646838272;
parameter    ap_ST_fsm_state79 = 85'd302231454903657293676544;
parameter    ap_ST_fsm_state80 = 85'd604462909807314587353088;
parameter    ap_ST_fsm_state81 = 85'd1208925819614629174706176;
parameter    ap_ST_fsm_state82 = 85'd2417851639229258349412352;
parameter    ap_ST_fsm_state83 = 85'd4835703278458516698824704;
parameter    ap_ST_fsm_state84 = 85'd9671406556917033397649408;
parameter    ap_ST_fsm_state85 = 85'd19342813113834066795298816;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [20:0] p_read;
input  [20:0] p_read1;
input  [20:0] p_read2;
output  [4:0] h_address0;
output   h_ce0;
input  [20:0] h_q0;
output  [4:0] h_address1;
output   h_ce1;
input  [20:0] h_q1;
output  [20:0] xk_admm_V_0;
output   xk_admm_V_0_ap_vld;

reg ap_idle;
reg[4:0] h_address0;
reg h_ce0;
reg[4:0] h_address1;
reg h_ce1;
reg xk_admm_V_0_ap_vld;

(* fsm_encoding = "none" *) reg   [84:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1_pp0_stage0_iter0;
wire   [0:0] icmp_ln74_fu_1292_p2;
reg    ap_condition_exit_pp0_iter0_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire    ap_CS_fsm_state85;
wire    ap_block_state85_pp0_stage84_iter0;
reg   [4:0] zk_admm_V_address0;
reg    zk_admm_V_ce0;
reg    zk_admm_V_we0;
reg   [20:0] zk_admm_V_d0;
wire   [20:0] zk_admm_V_q0;
reg   [4:0] zk_admm_V_address1;
reg    zk_admm_V_ce1;
reg    zk_admm_V_we1;
reg   [20:0] zk_admm_V_d1;
wire   [20:0] zk_admm_V_q1;
reg   [4:0] uk_admm_V_address0;
reg    uk_admm_V_ce0;
reg    uk_admm_V_we0;
reg   [20:0] uk_admm_V_d0;
wire   [20:0] uk_admm_V_q0;
reg   [4:0] uk_admm_V_address1;
reg    uk_admm_V_ce1;
reg    uk_admm_V_we1;
reg   [20:0] uk_admm_V_d1;
wire   [20:0] uk_admm_V_q1;
reg  signed [20:0] reg_1200;
wire    ap_CS_fsm_state2;
wire    ap_block_state2_pp0_stage1_iter0;
wire    ap_CS_fsm_state23;
wire    ap_block_state23_pp0_stage22_iter0;
reg  signed [20:0] reg_1204;
reg  signed [20:0] reg_1208;
wire    ap_CS_fsm_state3;
wire    ap_block_state3_pp0_stage2_iter0;
wire    ap_CS_fsm_state24;
wire    ap_block_state24_pp0_stage23_iter0;
reg  signed [20:0] reg_1212;
reg  signed [20:0] reg_1216;
wire    ap_CS_fsm_state4;
wire    ap_block_state4_pp0_stage3_iter0;
wire    ap_CS_fsm_state25;
wire    ap_block_state25_pp0_stage24_iter0;
reg  signed [20:0] reg_1220;
reg  signed [20:0] reg_1224;
wire    ap_CS_fsm_state5;
wire    ap_block_state5_pp0_stage4_iter0;
wire    ap_CS_fsm_state26;
wire    ap_block_state26_pp0_stage25_iter0;
reg  signed [20:0] reg_1228;
reg  signed [20:0] reg_1232;
wire    ap_CS_fsm_state6;
wire    ap_block_state6_pp0_stage5_iter0;
wire    ap_CS_fsm_state27;
wire    ap_block_state27_pp0_stage26_iter0;
reg  signed [20:0] reg_1236;
reg  signed [20:0] reg_1240;
wire    ap_CS_fsm_state7;
wire    ap_block_state7_pp0_stage6_iter0;
wire    ap_CS_fsm_state28;
wire    ap_block_state28_pp0_stage27_iter0;
reg  signed [20:0] reg_1244;
reg  signed [20:0] reg_1248;
wire    ap_CS_fsm_state8;
wire    ap_block_state8_pp0_stage7_iter0;
wire    ap_CS_fsm_state29;
wire    ap_block_state29_pp0_stage28_iter0;
reg  signed [20:0] reg_1252;
reg  signed [20:0] reg_1256;
wire    ap_CS_fsm_state9;
wire    ap_block_state9_pp0_stage8_iter0;
wire    ap_CS_fsm_state30;
wire    ap_block_state30_pp0_stage29_iter0;
reg  signed [20:0] reg_1260;
reg  signed [20:0] reg_1264;
wire    ap_CS_fsm_state10;
wire    ap_block_state10_pp0_stage9_iter0;
wire    ap_CS_fsm_state31;
wire    ap_block_state31_pp0_stage30_iter0;
reg  signed [20:0] reg_1268;
wire  signed [21:0] sext_ln813_71_fu_1272_p1;
reg  signed [21:0] sext_ln813_71_reg_21983;
wire  signed [21:0] sext_ln813_72_fu_1276_p1;
reg  signed [21:0] sext_ln813_72_reg_21988;
wire  signed [21:0] sext_ln813_73_fu_1280_p1;
reg  signed [21:0] sext_ln813_73_reg_21993;
wire    ap_CS_fsm_state13;
wire    ap_block_state13_pp0_stage12_iter0;
wire  signed [34:0] sext_ln1273_2_fu_1597_p1;
wire    ap_CS_fsm_state14;
wire    ap_block_state14_pp0_stage13_iter0;
wire  signed [34:0] sext_ln1273_6_fu_1601_p1;
wire  signed [20:0] select_ln302_3_fu_1671_p3;
reg  signed [20:0] select_ln302_3_reg_22388;
wire    ap_CS_fsm_state15;
wire    ap_block_state15_pp0_stage14_iter0;
wire  signed [20:0] select_ln302_5_fu_1741_p3;
reg  signed [20:0] select_ln302_5_reg_22394;
reg   [0:0] tmp_91_reg_22405;
reg   [0:0] tmp_183_reg_22420;
wire  signed [27:0] grp_fu_21397_p2;
reg  signed [27:0] mul_ln1273_1_reg_22425;
wire    ap_CS_fsm_state16;
wire    ap_block_state16_pp0_stage15_iter0;
wire   [20:0] select_ln346_36_fu_2155_p3;
reg   [20:0] select_ln346_36_reg_22431;
reg   [0:0] tmp_79_reg_22436;
wire  signed [20:0] select_ln302_9_fu_2310_p3;
reg  signed [20:0] select_ln302_9_reg_22451;
wire    ap_CS_fsm_state17;
wire    ap_block_state17_pp0_stage16_iter0;
wire  signed [34:0] grp_fu_21404_p2;
reg  signed [34:0] mul_ln1273_2_reg_22457;
wire   [20:0] select_ln346_38_fu_2522_p3;
reg   [20:0] select_ln346_38_reg_22463;
reg   [0:0] tmp_85_reg_22468;
wire  signed [33:0] grp_fu_21411_p2;
reg  signed [33:0] mul_ln1273_3_reg_22473;
reg   [0:0] tmp_97_reg_22479;
wire  signed [34:0] sext_ln1273_12_fu_2544_p1;
wire   [20:0] select_ln346_72_fu_2730_p3;
reg   [20:0] select_ln346_72_reg_22495;
wire  signed [34:0] grp_fu_21430_p2;
reg  signed [34:0] mul_ln1273_14_reg_22500;
reg   [0:0] tmp_177_reg_22506;
wire   [20:0] select_ln346_104_fu_2923_p3;
reg   [20:0] select_ln346_104_reg_22511;
wire  signed [20:0] select_ln302_11_fu_3063_p3;
reg  signed [20:0] select_ln302_11_reg_22516;
wire    ap_CS_fsm_state18;
wire    ap_block_state18_pp0_stage17_iter0;
wire   [20:0] select_ln346_40_fu_3271_p3;
reg   [20:0] select_ln346_40_reg_22522;
wire  signed [29:0] grp_fu_21449_p2;
reg  signed [29:0] mul_ln1273_4_reg_22527;
reg   [0:0] tmp_103_reg_22533;
wire  signed [34:0] sext_ln1273_16_fu_3286_p1;
wire   [0:0] tmp_169_fu_3331_p3;
reg   [0:0] tmp_169_reg_22559;
wire   [0:0] tmp_170_fu_3349_p3;
reg   [0:0] tmp_170_reg_22564;
wire   [20:0] add_ln377_15_fu_3368_p2;
reg   [20:0] add_ln377_15_reg_22569;
wire   [0:0] xor_ln896_34_fu_3382_p2;
reg   [0:0] xor_ln896_34_reg_22574;
wire   [0:0] tmp_173_fu_3388_p3;
reg   [0:0] tmp_173_reg_22579;
wire   [0:0] and_ln895_54_fu_3458_p2;
reg   [0:0] and_ln895_54_reg_22584;
wire   [0:0] or_ln896_15_fu_3470_p2;
reg   [0:0] or_ln896_15_reg_22590;
wire   [0:0] tmp_241_fu_3505_p3;
reg   [0:0] tmp_241_reg_22595;
wire   [0:0] tmp_242_fu_3523_p3;
reg   [0:0] tmp_242_reg_22600;
wire   [20:0] add_ln377_25_fu_3542_p2;
reg   [20:0] add_ln377_25_reg_22605;
wire   [0:0] xor_ln896_60_fu_3556_p2;
reg   [0:0] xor_ln896_60_reg_22610;
wire   [0:0] tmp_245_fu_3562_p3;
reg   [0:0] tmp_245_reg_22615;
wire   [0:0] and_ln895_70_fu_3632_p2;
reg   [0:0] and_ln895_70_reg_22620;
wire   [0:0] or_ln896_25_fu_3644_p2;
reg   [0:0] or_ln896_25_reg_22626;
wire   [20:0] add_ln377_3_fu_3878_p2;
reg   [20:0] add_ln377_3_reg_22631;
wire    ap_CS_fsm_state19;
wire    ap_block_state19_pp0_stage18_iter0;
wire   [0:0] and_ln895_38_fu_3980_p2;
reg   [0:0] and_ln895_38_reg_22636;
wire   [0:0] or_ln346_3_fu_4010_p2;
reg   [0:0] or_ln346_3_reg_22641;
wire  signed [34:0] grp_fu_21474_p2;
reg  signed [34:0] mul_ln1273_5_reg_22646;
reg   [0:0] tmp_109_reg_22652;
wire  signed [27:0] grp_fu_21481_p2;
reg  signed [27:0] mul_ln1273_6_reg_22657;
reg   [0:0] tmp_115_reg_22663;
wire   [20:0] add_ln377_16_fu_4127_p2;
reg   [20:0] add_ln377_16_reg_22673;
wire   [0:0] and_ln895_55_fu_4229_p2;
reg   [0:0] and_ln895_55_reg_22678;
wire   [0:0] or_ln346_16_fu_4259_p2;
reg   [0:0] or_ln346_16_reg_22683;
wire   [20:0] select_ln346_114_fu_4499_p3;
reg   [20:0] select_ln346_114_reg_22693;
wire   [20:0] select_ln346_44_fu_4865_p3;
reg   [20:0] select_ln346_44_reg_22698;
wire    ap_CS_fsm_state20;
wire    ap_block_state20_pp0_stage19_iter0;
wire  signed [34:0] grp_fu_21488_p2;
reg  signed [34:0] mul_ln1273_7_reg_22703;
reg   [0:0] tmp_121_reg_22709;
wire   [20:0] add_ln377_17_fu_4986_p2;
reg   [20:0] add_ln377_17_reg_22719;
wire   [0:0] and_ln895_56_fu_5088_p2;
reg   [0:0] and_ln895_56_reg_22724;
wire   [0:0] or_ln346_17_fu_5118_p2;
reg   [0:0] or_ln346_17_reg_22729;
wire  signed [34:0] grp_fu_21495_p2;
reg  signed [34:0] mul_ln1273_15_reg_22734;
reg   [0:0] tmp_193_reg_22740;
wire  signed [27:0] grp_fu_21502_p2;
reg  signed [27:0] mul_ln1273_16_reg_22745;
reg   [0:0] tmp_199_reg_22751;
wire   [20:0] select_ln346_46_fu_5486_p3;
reg   [20:0] select_ln346_46_reg_22761;
wire    ap_CS_fsm_state21;
wire    ap_block_state21_pp0_stage20_iter0;
wire  signed [33:0] grp_fu_21509_p2;
reg  signed [33:0] mul_ln1273_8_reg_22766;
reg   [0:0] tmp_133_reg_22772;
wire  signed [29:0] grp_fu_21516_p2;
reg  signed [29:0] mul_ln1273_9_reg_22777;
reg   [0:0] tmp_139_reg_22783;
wire   [0:0] tmp_191_fu_5647_p3;
reg   [0:0] tmp_191_reg_22788;
wire   [0:0] tmp_192_fu_5665_p3;
reg   [0:0] tmp_192_reg_22793;
wire   [20:0] add_ln377_18_fu_5676_p2;
reg   [20:0] add_ln377_18_reg_22798;
wire   [0:0] xor_ln896_42_fu_5690_p2;
reg   [0:0] xor_ln896_42_reg_22803;
wire   [0:0] tmp_195_fu_5696_p3;
reg   [0:0] tmp_195_reg_22808;
wire   [0:0] and_ln895_59_fu_5766_p2;
reg   [0:0] and_ln895_59_reg_22813;
wire   [0:0] or_ln896_18_fu_5778_p2;
reg   [0:0] or_ln896_18_reg_22819;
wire  signed [34:0] grp_fu_21523_p2;
reg  signed [34:0] mul_ln1273_17_reg_22824;
reg   [0:0] tmp_205_reg_22830;
wire   [0:0] tmp_255_fu_5820_p3;
reg   [0:0] tmp_255_reg_22840;
wire   [0:0] tmp_256_fu_5838_p3;
reg   [0:0] tmp_256_reg_22845;
wire   [20:0] add_ln377_26_fu_5857_p2;
reg   [20:0] add_ln377_26_reg_22850;
wire   [0:0] xor_ln896_66_fu_5871_p2;
reg   [0:0] xor_ln896_66_reg_22855;
wire   [0:0] tmp_259_fu_5877_p3;
reg   [0:0] tmp_259_reg_22860;
wire   [0:0] and_ln895_75_fu_5947_p2;
reg   [0:0] and_ln895_75_reg_22865;
wire   [0:0] or_ln896_26_fu_5959_p2;
reg   [0:0] or_ln896_26_reg_22871;
wire  signed [27:0] grp_fu_21539_p2;
reg  signed [27:0] mul_ln1273_23_reg_22876;
reg   [0:0] tmp_263_reg_22882;
wire   [20:0] select_ln346_48_fu_6176_p3;
reg   [20:0] select_ln346_48_reg_22892;
wire    ap_CS_fsm_state22;
wire    ap_block_state22_pp0_stage21_iter0;
wire  signed [35:0] grp_fu_21546_p2;
reg  signed [35:0] mul_ln1273_10_reg_22897;
reg   [0:0] tmp_145_reg_22902;
wire   [20:0] add_ln377_19_fu_6288_p2;
reg   [20:0] add_ln377_19_reg_22907;
wire   [0:0] and_ln895_60_fu_6390_p2;
reg   [0:0] and_ln895_60_reg_22912;
wire   [0:0] or_ln346_19_fu_6420_p2;
reg   [0:0] or_ln346_19_reg_22917;
wire  signed [35:0] grp_fu_21553_p2;
reg  signed [35:0] mul_ln1273_18_reg_22922;
reg   [0:0] tmp_219_reg_22927;
wire   [20:0] add_ln377_27_fu_6530_p2;
reg   [20:0] add_ln377_27_reg_22932;
wire   [0:0] and_ln895_76_fu_6632_p2;
reg   [0:0] and_ln895_76_reg_22937;
wire   [0:0] or_ln346_27_fu_6662_p2;
reg   [0:0] or_ln346_27_reg_22942;
wire   [20:0] select_ln346_50_fu_6872_p3;
reg   [20:0] select_ln346_50_reg_22947;
wire  signed [35:0] grp_fu_21560_p2;
reg  signed [35:0] mul_ln1273_11_reg_22952;
reg   [0:0] tmp_155_reg_22957;
wire   [20:0] select_ln346_88_fu_7101_p3;
reg   [20:0] select_ln346_88_reg_22962;
wire   [0:0] tmp_271_fu_7239_p3;
reg   [0:0] tmp_271_reg_22967;
wire   [0:0] tmp_272_fu_7257_p3;
reg   [0:0] tmp_272_reg_22972;
wire   [20:0] add_ln377_28_fu_7276_p2;
reg   [20:0] add_ln377_28_reg_22977;
wire   [0:0] xor_ln896_72_fu_7290_p2;
reg   [0:0] xor_ln896_72_reg_22982;
wire   [0:0] tmp_275_fu_7296_p3;
reg   [0:0] tmp_275_reg_22987;
wire   [0:0] and_ln895_79_fu_7366_p2;
reg   [0:0] and_ln895_79_reg_22992;
wire   [0:0] or_ln896_28_fu_7378_p2;
reg   [0:0] or_ln896_28_reg_22998;
wire   [20:0] select_ln346_52_fu_7584_p3;
reg   [20:0] select_ln346_52_reg_23003;
wire   [20:0] add_ln377_21_fu_7689_p2;
reg   [20:0] add_ln377_21_reg_23008;
wire   [0:0] and_ln895_62_fu_7791_p2;
reg   [0:0] and_ln895_62_reg_23013;
wire   [0:0] or_ln346_21_fu_7821_p2;
reg   [0:0] or_ln346_21_reg_23018;
wire  signed [35:0] grp_fu_21575_p2;
reg  signed [35:0] mul_ln1273_19_reg_23023;
reg   [0:0] tmp_229_reg_23028;
wire   [0:0] tmp_281_fu_7989_p3;
reg   [0:0] tmp_281_reg_23033;
wire   [0:0] tmp_282_fu_8007_p3;
reg   [0:0] tmp_282_reg_23038;
wire   [20:0] add_ln377_29_fu_8026_p2;
reg   [20:0] add_ln377_29_reg_23043;
wire   [0:0] xor_ln896_76_fu_8040_p2;
reg   [0:0] xor_ln896_76_reg_23048;
wire   [0:0] tmp_285_fu_8046_p3;
reg   [0:0] tmp_285_reg_23053;
wire   [0:0] and_ln895_82_fu_8116_p2;
reg   [0:0] and_ln895_82_reg_23058;
wire   [0:0] or_ln896_29_fu_8128_p2;
reg   [0:0] or_ln896_29_reg_23064;
wire   [20:0] add_ln377_9_fu_8231_p2;
reg   [20:0] add_ln377_9_reg_23069;
wire   [0:0] and_ln895_44_fu_8333_p2;
reg   [0:0] and_ln895_44_reg_23074;
wire   [0:0] or_ln346_9_fu_8363_p2;
reg   [0:0] or_ln346_9_reg_23079;
wire   [20:0] add_ln377_22_fu_8478_p2;
reg   [20:0] add_ln377_22_reg_23084;
wire   [0:0] and_ln895_64_fu_8580_p2;
reg   [0:0] and_ln895_64_reg_23089;
wire   [0:0] or_ln346_22_fu_8610_p2;
reg   [0:0] or_ln346_22_reg_23094;
wire  signed [29:0] sext_ln1273_37_fu_8721_p1;
wire  signed [29:0] sub_ln1273_4_fu_8753_p2;
reg  signed [29:0] sub_ln1273_4_reg_23109;
reg   [0:0] tmp_325_reg_23115;
wire   [20:0] select_ln346_56_fu_8991_p3;
reg   [20:0] select_ln346_56_reg_23120;
wire   [20:0] add_ln377_23_fu_9158_p2;
reg   [20:0] add_ln377_23_reg_23125;
wire   [0:0] and_ln895_67_fu_9260_p2;
reg   [0:0] and_ln895_67_reg_23130;
wire   [0:0] or_ln346_23_fu_9290_p2;
reg   [0:0] or_ln346_23_reg_23135;
wire   [20:0] add_ln377_11_fu_9354_p2;
reg   [20:0] add_ln377_11_reg_23140;
wire   [0:0] and_ln895_46_fu_9456_p2;
reg   [0:0] and_ln895_46_reg_23145;
wire   [0:0] or_ln346_11_fu_9486_p2;
reg   [0:0] or_ln346_11_reg_23150;
wire  signed [20:0] select_ln302_22_fu_9610_p3;
reg  signed [20:0] select_ln302_22_reg_23155;
reg   [0:0] tmp_337_reg_23171;
wire   [20:0] add_ln377_12_fu_9715_p2;
reg   [20:0] add_ln377_12_reg_23176;
wire   [0:0] and_ln895_47_fu_9817_p2;
reg   [0:0] and_ln895_47_reg_23181;
wire   [0:0] or_ln346_12_fu_9847_p2;
reg   [0:0] or_ln346_12_reg_23186;
wire  signed [29:0] grp_fu_21590_p2;
reg  signed [29:0] mul_ln1273_28_reg_23191;
reg   [0:0] tmp_307_reg_23197;
wire  signed [34:0] grp_fu_21597_p2;
reg  signed [34:0] mul_ln1273_32_reg_23202;
reg   [0:0] tmp_343_reg_23208;
wire   [20:0] add_ln377_13_fu_10026_p2;
reg   [20:0] add_ln377_13_reg_23213;
wire   [0:0] and_ln895_50_fu_10128_p2;
reg   [0:0] and_ln895_50_reg_23218;
wire   [0:0] or_ln346_13_fu_10158_p2;
reg   [0:0] or_ln346_13_reg_23223;
wire  signed [30:0] grp_fu_21604_p2;
reg  signed [30:0] mul_ln1273_27_reg_23243;
reg   [0:0] tmp_301_reg_23249;
wire  signed [33:0] grp_fu_21611_p2;
reg  signed [33:0] mul_ln1273_30_reg_23254;
reg   [0:0] tmp_319_reg_23260;
wire   [20:0] select_ln346_135_fu_10548_p3;
reg   [20:0] select_ln346_135_reg_23265;
wire    ap_CS_fsm_state33;
wire    ap_block_state33_pp0_stage32_iter0;
wire  signed [17:0] add_ln377_33_fu_10594_p2;
reg  signed [17:0] add_ln377_33_reg_23270;
wire   [0:0] and_ln895_89_fu_10694_p2;
reg   [0:0] and_ln895_89_reg_23275;
wire   [0:0] or_ln346_33_fu_10724_p2;
reg   [0:0] or_ln346_33_reg_23280;
wire  signed [16:0] add_ln377_36_fu_10768_p2;
reg  signed [16:0] add_ln377_36_reg_23285;
wire   [0:0] and_ln895_92_fu_10868_p2;
reg   [0:0] and_ln895_92_reg_23290;
wire   [0:0] or_ln346_36_fu_10898_p2;
reg   [0:0] or_ln346_36_reg_23295;
wire   [20:0] select_ln346_137_fu_11111_p3;
reg   [20:0] select_ln346_137_reg_23300;
wire    ap_CS_fsm_state34;
wire    ap_block_state34_pp0_stage33_iter0;
wire   [20:0] select_ln346_143_fu_11341_p3;
reg   [20:0] select_ln346_143_reg_23305;
wire   [20:0] add_ln377_37_fu_11444_p2;
reg   [20:0] add_ln377_37_reg_23310;
wire   [0:0] and_ln895_93_fu_11546_p2;
reg   [0:0] and_ln895_93_reg_23315;
wire   [0:0] or_ln346_37_fu_11576_p2;
reg   [0:0] or_ln346_37_reg_23320;
wire   [20:0] add_ln377_32_fu_11640_p2;
reg   [20:0] add_ln377_32_reg_23325;
wire    ap_CS_fsm_state35;
wire    ap_block_state35_pp0_stage34_iter0;
wire   [0:0] and_ln895_88_fu_11742_p2;
reg   [0:0] and_ln895_88_reg_23330;
wire   [0:0] or_ln346_32_fu_11772_p2;
reg   [0:0] or_ln346_32_reg_23335;
wire   [20:0] add_ln377_35_fu_11836_p2;
reg   [20:0] add_ln377_35_reg_23340;
wire   [0:0] and_ln895_91_fu_11938_p2;
reg   [0:0] and_ln895_91_reg_23345;
wire   [0:0] or_ln346_35_fu_11968_p2;
reg   [0:0] or_ln346_35_reg_23350;
wire   [20:0] add_ln377_38_fu_12042_p2;
reg   [20:0] add_ln377_38_reg_23355;
wire   [0:0] and_ln895_94_fu_12144_p2;
reg   [0:0] and_ln895_94_reg_23360;
wire   [0:0] or_ln346_38_fu_12174_p2;
reg   [0:0] or_ln346_38_reg_23365;
wire  signed [20:0] select_ln346_139_fu_12187_p3;
reg  signed [20:0] select_ln346_139_reg_23370;
wire    ap_CS_fsm_state36;
wire    ap_block_state36_pp0_stage35_iter0;
wire  signed [20:0] select_ln346_145_fu_12206_p3;
reg  signed [20:0] select_ln346_145_reg_23375;
wire  signed [29:0] sext_ln1273_40_fu_12212_p1;
wire  signed [33:0] sext_ln1273_41_fu_12216_p1;
wire  signed [28:0] sext_ln1273_42_fu_12220_p1;
wire  signed [27:0] sext_ln1273_43_fu_12224_p1;
reg  signed [27:0] sext_ln1273_43_reg_23399;
wire  signed [34:0] sext_ln1273_44_fu_12228_p1;
reg  signed [34:0] sext_ln1273_44_reg_23405;
wire  signed [28:0] sext_ln1273_45_fu_12232_p1;
wire  signed [34:0] sext_ln1273_47_fu_12236_p1;
reg  signed [34:0] sext_ln1273_47_reg_23419;
wire  signed [20:0] select_ln346_151_fu_12531_p3;
reg  signed [20:0] select_ln346_151_reg_23427;
wire    ap_CS_fsm_state37;
wire    ap_block_state37_pp0_stage36_iter0;
wire  signed [27:0] sext_ln1273_46_fu_12537_p1;
wire  signed [27:0] sext_ln1273_48_fu_12540_p1;
wire  signed [34:0] sext_ln1273_49_fu_12544_p1;
wire   [20:0] add_ln377_39_fu_13145_p2;
reg   [20:0] add_ln377_39_reg_23450;
wire    ap_CS_fsm_state39;
wire    ap_block_state39_pp0_stage38_iter0;
wire   [0:0] and_ln895_95_fu_13245_p2;
reg   [0:0] and_ln895_95_reg_23455;
wire   [0:0] or_ln346_39_fu_13275_p2;
reg   [0:0] or_ln346_39_reg_23460;
wire  signed [14:0] add_ln377_40_fu_13319_p2;
reg  signed [14:0] add_ln377_40_reg_23465;
wire   [0:0] and_ln895_98_fu_13419_p2;
reg   [0:0] and_ln895_98_reg_23470;
wire   [0:0] or_ln346_40_fu_13449_p2;
reg   [0:0] or_ln346_40_reg_23475;
wire   [20:0] select_ln346_165_fu_13633_p3;
reg   [20:0] select_ln346_165_reg_23480;
wire  signed [15:0] add_ln377_43_fu_13679_p2;
reg  signed [15:0] add_ln377_43_reg_23485;
wire   [0:0] and_ln895_104_fu_13779_p2;
reg   [0:0] and_ln895_104_reg_23490;
wire   [0:0] or_ln346_43_fu_13809_p2;
reg   [0:0] or_ln346_43_reg_23495;
wire  signed [34:0] grp_fu_21714_p2;
reg  signed [34:0] mul_ln1273_40_reg_23500;
wire   [20:0] select_ln346_177_fu_13997_p3;
reg   [20:0] select_ln346_177_reg_23506;
reg   [0:0] tmp_403_reg_23511;
wire  signed [16:0] add_ln377_48_fu_14050_p2;
reg  signed [16:0] add_ln377_48_reg_23516;
wire   [0:0] and_ln895_110_fu_14150_p2;
reg   [0:0] and_ln895_110_reg_23521;
wire   [0:0] or_ln346_48_fu_14180_p2;
reg   [0:0] or_ln346_48_reg_23526;
wire  signed [28:0] grp_fu_21733_p2;
reg  signed [28:0] mul_ln1273_43_reg_23531;
reg   [0:0] tmp_421_reg_23537;
wire   [20:0] select_ln346_201_fu_14371_p3;
reg   [20:0] select_ln346_201_reg_23542;
wire  signed [15:0] add_ln377_55_fu_14417_p2;
reg  signed [15:0] add_ln377_55_reg_23547;
wire   [0:0] and_ln895_122_fu_14517_p2;
reg   [0:0] and_ln895_122_reg_23552;
wire   [0:0] or_ln346_55_fu_14547_p2;
reg   [0:0] or_ln346_55_reg_23557;
wire  signed [34:0] grp_fu_21776_p2;
reg  signed [34:0] mul_ln1273_52_reg_23562;
wire   [20:0] select_ln346_213_fu_14735_p3;
reg   [20:0] select_ln346_213_reg_23568;
reg   [0:0] tmp_487_reg_23573;
wire  signed [16:0] add_ln377_60_fu_14788_p2;
reg  signed [16:0] add_ln377_60_reg_23578;
wire   [0:0] and_ln895_128_fu_14888_p2;
reg   [0:0] and_ln895_128_reg_23583;
wire   [0:0] or_ln346_60_fu_14918_p2;
reg   [0:0] or_ln346_60_reg_23588;
wire  signed [28:0] grp_fu_21795_p2;
reg  signed [28:0] mul_ln1273_55_reg_23593;
reg   [0:0] tmp_505_reg_23599;
wire   [0:0] tmp_373_fu_15188_p3;
reg   [0:0] tmp_373_reg_23604;
wire    ap_CS_fsm_state40;
wire    ap_block_state40_pp0_stage39_iter0;
wire   [0:0] tmp_374_fu_15206_p3;
reg   [0:0] tmp_374_reg_23609;
wire   [20:0] add_ln377_42_fu_15225_p2;
reg   [20:0] add_ln377_42_reg_23614;
wire   [0:0] xor_ln896_106_fu_15239_p2;
reg   [0:0] xor_ln896_106_reg_23619;
wire   [0:0] tmp_377_fu_15245_p3;
reg   [0:0] tmp_377_reg_23624;
wire   [0:0] and_ln895_102_fu_15315_p2;
reg   [0:0] and_ln895_102_reg_23629;
wire   [0:0] or_ln896_42_fu_15327_p2;
reg   [0:0] or_ln896_42_reg_23635;
wire   [0:0] tmp_387_fu_15380_p3;
reg   [0:0] tmp_387_reg_23640;
wire   [0:0] tmp_388_fu_15398_p3;
reg   [0:0] tmp_388_reg_23645;
wire   [20:0] add_ln377_44_fu_15417_p2;
reg   [20:0] add_ln377_44_reg_23650;
wire   [0:0] xor_ln896_111_fu_15431_p2;
reg   [0:0] xor_ln896_111_reg_23655;
wire   [0:0] tmp_391_fu_15437_p3;
reg   [0:0] tmp_391_reg_23660;
wire   [0:0] and_ln895_105_fu_15507_p2;
reg   [0:0] and_ln895_105_reg_23665;
wire   [0:0] or_ln896_44_fu_15519_p2;
reg   [0:0] or_ln896_44_reg_23671;
wire  signed [34:0] grp_fu_21819_p2;
reg  signed [34:0] mul_ln1273_41_reg_23676;
wire   [20:0] select_ln346_179_fu_15725_p3;
reg   [20:0] select_ln346_179_reg_23682;
reg   [0:0] tmp_409_reg_23687;
wire  signed [27:0] grp_fu_21826_p2;
reg  signed [27:0] mul_ln1273_44_reg_23692;
wire   [20:0] select_ln346_185_fu_15962_p3;
reg   [20:0] select_ln346_185_reg_23698;
reg   [0:0] tmp_427_reg_23703;
wire   [20:0] add_ln377_51_fu_16011_p2;
reg   [20:0] add_ln377_51_reg_23708;
wire   [0:0] and_ln895_113_fu_16111_p2;
reg   [0:0] and_ln895_113_reg_23713;
wire   [0:0] or_ln346_51_fu_16141_p2;
reg   [0:0] or_ln346_51_reg_23718;
wire  signed [14:0] add_ln377_52_fu_16185_p2;
reg  signed [14:0] add_ln377_52_reg_23723;
wire   [0:0] and_ln895_116_fu_16285_p2;
reg   [0:0] and_ln895_116_reg_23728;
wire   [0:0] or_ln346_52_fu_16315_p2;
reg   [0:0] or_ln346_52_reg_23733;
wire   [0:0] tmp_457_fu_16346_p3;
reg   [0:0] tmp_457_reg_23738;
wire   [0:0] tmp_458_fu_16364_p3;
reg   [0:0] tmp_458_reg_23743;
wire   [20:0] add_ln377_54_fu_16383_p2;
reg   [20:0] add_ln377_54_reg_23748;
wire   [0:0] xor_ln896_136_fu_16397_p2;
reg   [0:0] xor_ln896_136_reg_23753;
wire   [0:0] tmp_461_fu_16403_p3;
reg   [0:0] tmp_461_reg_23758;
wire   [0:0] and_ln895_120_fu_16473_p2;
reg   [0:0] and_ln895_120_reg_23763;
wire   [0:0] or_ln896_54_fu_16485_p2;
reg   [0:0] or_ln896_54_reg_23769;
wire   [0:0] tmp_471_fu_16538_p3;
reg   [0:0] tmp_471_reg_23774;
wire   [0:0] tmp_472_fu_16556_p3;
reg   [0:0] tmp_472_reg_23779;
wire   [20:0] add_ln377_56_fu_16575_p2;
reg   [20:0] add_ln377_56_reg_23784;
wire   [0:0] xor_ln896_141_fu_16589_p2;
reg   [0:0] xor_ln896_141_reg_23789;
wire   [0:0] tmp_475_fu_16595_p3;
reg   [0:0] tmp_475_reg_23794;
wire   [0:0] and_ln895_123_fu_16665_p2;
reg   [0:0] and_ln895_123_reg_23799;
wire   [0:0] or_ln896_56_fu_16677_p2;
reg   [0:0] or_ln896_56_reg_23805;
wire  signed [34:0] grp_fu_21872_p2;
reg  signed [34:0] mul_ln1273_53_reg_23810;
wire   [20:0] select_ln346_215_fu_16883_p3;
reg   [20:0] select_ln346_215_reg_23816;
reg   [0:0] tmp_493_reg_23821;
wire  signed [27:0] grp_fu_21879_p2;
reg  signed [27:0] mul_ln1273_56_reg_23826;
wire   [20:0] select_ln346_221_fu_17120_p3;
reg   [20:0] select_ln346_221_reg_23832;
reg   [0:0] tmp_511_reg_23837;
wire   [20:0] select_ln346_169_fu_17215_p3;
reg   [20:0] select_ln346_169_reg_23842;
wire    ap_CS_fsm_state41;
wire    ap_block_state41_pp0_stage40_iter0;
wire   [20:0] select_ln346_175_fu_17303_p3;
reg   [20:0] select_ln346_175_reg_23847;
wire   [20:0] select_ln346_181_fu_17511_p3;
reg   [20:0] select_ln346_181_reg_23852;
wire   [20:0] select_ln346_187_fu_17723_p3;
reg   [20:0] select_ln346_187_reg_23857;
wire   [20:0] select_ln346_205_fu_18043_p3;
reg   [20:0] select_ln346_205_reg_23862;
wire   [20:0] select_ln346_211_fu_18131_p3;
reg   [20:0] select_ln346_211_reg_23867;
wire   [20:0] select_ln346_217_fu_18339_p3;
reg   [20:0] select_ln346_217_reg_23872;
wire   [20:0] select_ln346_223_fu_18551_p3;
reg   [20:0] select_ln346_223_reg_23877;
reg  signed [20:0] zk_admm_V_load_reg_23882;
wire    ap_CS_fsm_state67;
wire    ap_block_state67_pp0_stage66_iter0;
reg  signed [20:0] zk_admm_V_load_1_reg_23888;
reg  signed [20:0] zk_admm_V_load_2_reg_23894;
wire    ap_CS_fsm_state68;
wire    ap_block_state68_pp0_stage67_iter0;
reg  signed [20:0] zk_admm_V_load_3_reg_23900;
reg  signed [20:0] zk_admm_V_load_4_reg_23906;
wire    ap_CS_fsm_state69;
wire    ap_block_state69_pp0_stage68_iter0;
reg  signed [20:0] zk_admm_V_load_5_reg_23912;
reg  signed [20:0] zk_admm_V_load_6_reg_23918;
wire    ap_CS_fsm_state70;
wire    ap_block_state70_pp0_stage69_iter0;
reg  signed [20:0] zk_admm_V_load_7_reg_23924;
reg  signed [20:0] zk_admm_V_load_8_reg_23930;
wire    ap_CS_fsm_state71;
wire    ap_block_state71_pp0_stage70_iter0;
reg  signed [20:0] zk_admm_V_load_9_reg_23936;
reg  signed [20:0] zk_admm_V_load_10_reg_23942;
wire    ap_CS_fsm_state72;
wire    ap_block_state72_pp0_stage71_iter0;
reg  signed [20:0] zk_admm_V_load_11_reg_23948;
reg  signed [20:0] zk_admm_V_load_12_reg_23954;
wire    ap_CS_fsm_state73;
wire    ap_block_state73_pp0_stage72_iter0;
reg  signed [20:0] zk_admm_V_load_13_reg_23960;
reg  signed [20:0] zk_admm_V_load_14_reg_23966;
wire    ap_CS_fsm_state74;
wire    ap_block_state74_pp0_stage73_iter0;
reg  signed [20:0] zk_admm_V_load_15_reg_23972;
reg  signed [20:0] zk_admm_V_load_16_reg_23978;
wire    ap_CS_fsm_state75;
wire    ap_block_state75_pp0_stage74_iter0;
reg  signed [20:0] zk_admm_V_load_17_reg_23984;
reg   [4:0] temp_address0;
reg    temp_ce0;
reg    temp_we0;
wire   [20:0] temp_q0;
reg   [4:0] temp_address1;
reg    temp_ce1;
reg    temp_we1;
wire   [20:0] temp_q1;
reg   [4:0] Hxk_V_address0;
reg    Hxk_V_ce0;
reg    Hxk_V_we0;
reg   [20:0] Hxk_V_d0;
wire   [20:0] Hxk_V_q0;
reg   [4:0] Hxk_V_address1;
reg    Hxk_V_ce1;
reg    Hxk_V_we1;
reg   [20:0] Hxk_V_d1;
wire   [20:0] Hxk_V_q1;
reg   [4:0] temp4_V_address0;
reg    temp4_V_ce0;
reg    temp4_V_we0;
wire   [20:0] temp4_V_q0;
reg   [4:0] temp4_V_address1;
reg    temp4_V_ce1;
reg    temp4_V_we1;
wire   [20:0] temp4_V_q1;
reg   [4:0] temp5_address0;
reg    temp5_ce0;
reg    temp5_we0;
wire   [20:0] temp5_q0;
reg   [4:0] temp5_address1;
reg    temp5_ce1;
reg    temp5_we1;
wire   [20:0] temp5_q1;
reg   [4:0] temp6_V_address0;
reg    temp6_V_ce0;
reg    temp6_V_we0;
reg   [20:0] temp6_V_d0;
wire   [20:0] temp6_V_q0;
reg   [4:0] temp6_V_address1;
reg    temp6_V_ce1;
reg    temp6_V_we1;
reg   [20:0] temp6_V_d1;
wire   [20:0] temp6_V_q1;
reg   [4:0] temp7_address0;
reg    temp7_ce0;
reg    temp7_we0;
wire   [20:0] temp7_q0;
reg   [4:0] temp7_address1;
reg    temp7_ce1;
reg    temp7_we1;
wire   [20:0] temp7_q1;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_done;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_idle;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_ready;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0;
reg   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1;
reg   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address0;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce0;
reg   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address1;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce1;
reg   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0;
wire   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0;
wire   [4:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1;
wire    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1;
wire   [20:0] grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1;
reg    grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg;
reg   [84:0] ap_NS_fsm;
wire    ap_NS_fsm_state2;
wire    ap_CS_fsm_state11;
wire    ap_NS_fsm_state12;
wire    ap_CS_fsm_state45;
wire    ap_NS_fsm_state46;
wire    ap_CS_fsm_state65;
wire    ap_NS_fsm_state66;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state46;
wire    ap_CS_fsm_state47;
wire    ap_CS_fsm_state48;
wire    ap_CS_fsm_state49;
wire    ap_CS_fsm_state50;
wire    ap_CS_fsm_state51;
wire    ap_CS_fsm_state52;
wire    ap_CS_fsm_state53;
wire    ap_CS_fsm_state54;
wire    ap_CS_fsm_state55;
wire    ap_CS_fsm_state66;
reg   [4:0] i_fu_310;
wire   [4:0] i_2_fu_1298_p2;
wire    ap_loop_init;
reg   [4:0] ap_sig_allocacmp_i_1;
wire    ap_CS_fsm_state77;
wire    ap_block_state77_pp0_stage76_iter0;
wire   [20:0] select_ln302_42_fu_20203_p3;
wire   [20:0] select_ln302_43_fu_20272_p3;
wire    ap_CS_fsm_state78;
wire    ap_block_state78_pp0_stage77_iter0;
wire   [20:0] select_ln302_44_fu_20341_p3;
wire   [20:0] select_ln302_45_fu_20410_p3;
wire    ap_CS_fsm_state79;
wire    ap_block_state79_pp0_stage78_iter0;
wire   [20:0] select_ln302_46_fu_20479_p3;
wire   [20:0] select_ln302_47_fu_20548_p3;
wire    ap_CS_fsm_state80;
wire    ap_block_state80_pp0_stage79_iter0;
wire   [20:0] select_ln302_48_fu_20617_p3;
wire   [20:0] select_ln302_49_fu_20686_p3;
wire    ap_CS_fsm_state81;
wire    ap_block_state81_pp0_stage80_iter0;
wire   [20:0] select_ln302_50_fu_20755_p3;
wire   [20:0] select_ln302_51_fu_20824_p3;
wire    ap_CS_fsm_state82;
wire    ap_block_state82_pp0_stage81_iter0;
wire   [20:0] select_ln302_52_fu_20893_p3;
wire   [20:0] select_ln302_53_fu_20962_p3;
wire    ap_CS_fsm_state83;
wire    ap_block_state83_pp0_stage82_iter0;
wire   [20:0] select_ln302_54_fu_21031_p3;
wire   [20:0] select_ln302_55_fu_21100_p3;
wire    ap_CS_fsm_state84;
wire    ap_block_state84_pp0_stage83_iter0;
wire   [20:0] select_ln302_56_fu_21169_p3;
wire   [20:0] select_ln302_57_fu_21238_p3;
wire   [20:0] select_ln302_58_fu_21307_p3;
wire   [20:0] select_ln302_59_fu_21376_p3;
wire    ap_block_state12_pp0_stage11_iter0;
wire   [20:0] select_ln346_229_fu_12382_p3;
wire   [20:0] select_ln346_233_fu_12515_p3;
wire   [20:0] select_ln346_235_fu_12622_p3;
wire   [20:0] select_ln346_241_fu_12832_p3;
wire    ap_CS_fsm_state38;
wire    ap_block_state38_pp0_stage37_iter0;
wire   [20:0] select_ln346_245_fu_13003_p3;
wire   [20:0] select_ln346_247_fu_13102_p3;
wire   [20:0] select_ln346_157_fu_15036_p3;
wire   [20:0] select_ln346_163_fu_15154_p3;
wire   [20:0] select_ln346_193_fu_17836_p3;
wire   [20:0] select_ln346_199_fu_17954_p3;
wire    ap_CS_fsm_state42;
wire    ap_block_state42_pp0_stage41_iter0;
wire    ap_CS_fsm_state43;
wire    ap_block_state43_pp0_stage42_iter0;
wire    ap_CS_fsm_state44;
wire    ap_block_state44_pp0_stage43_iter0;
wire    ap_block_state45_pp0_stage44_iter0;
wire    ap_CS_fsm_state56;
wire    ap_block_state56_pp0_stage55_iter0;
wire    ap_CS_fsm_state57;
wire    ap_block_state57_pp0_stage56_iter0;
wire    ap_CS_fsm_state58;
wire    ap_block_state58_pp0_stage57_iter0;
wire    ap_CS_fsm_state59;
wire    ap_block_state59_pp0_stage58_iter0;
wire    ap_CS_fsm_state60;
wire    ap_block_state60_pp0_stage59_iter0;
wire    ap_CS_fsm_state61;
wire    ap_block_state61_pp0_stage60_iter0;
wire    ap_CS_fsm_state62;
wire    ap_block_state62_pp0_stage61_iter0;
wire    ap_CS_fsm_state63;
wire    ap_block_state63_pp0_stage62_iter0;
wire    ap_CS_fsm_state64;
wire    ap_block_state64_pp0_stage63_iter0;
wire   [20:0] select_ln302_24_fu_18621_p3;
wire   [20:0] select_ln302_25_fu_18692_p3;
wire   [20:0] select_ln302_26_fu_18797_p3;
wire   [20:0] select_ln302_27_fu_18868_p3;
wire   [20:0] select_ln302_28_fu_18973_p3;
wire   [20:0] select_ln302_29_fu_19044_p3;
wire   [20:0] select_ln302_30_fu_19149_p3;
wire   [20:0] select_ln302_31_fu_19220_p3;
wire   [20:0] select_ln302_32_fu_19325_p3;
wire   [20:0] select_ln302_33_fu_19396_p3;
wire   [20:0] select_ln302_34_fu_19501_p3;
wire   [20:0] select_ln302_35_fu_19572_p3;
wire   [20:0] select_ln302_36_fu_19677_p3;
wire   [20:0] select_ln302_37_fu_19748_p3;
wire   [20:0] select_ln302_38_fu_19853_p3;
wire   [20:0] select_ln302_39_fu_19924_p3;
wire    ap_block_state65_pp0_stage64_iter0;
wire   [20:0] select_ln302_40_fu_20029_p3;
wire   [20:0] select_ln302_41_fu_20100_p3;
wire   [20:0] zext_ln50_fu_18713_p1;
wire   [20:0] zext_ln50_1_fu_18730_p1;
wire   [20:0] zext_ln50_2_fu_18889_p1;
wire   [20:0] zext_ln50_3_fu_18906_p1;
wire   [20:0] zext_ln50_4_fu_19065_p1;
wire   [20:0] zext_ln50_5_fu_19082_p1;
wire   [20:0] zext_ln50_6_fu_19241_p1;
wire   [20:0] zext_ln50_7_fu_19258_p1;
wire   [20:0] zext_ln50_8_fu_19417_p1;
wire   [20:0] zext_ln50_9_fu_19434_p1;
wire   [20:0] zext_ln50_10_fu_19593_p1;
wire   [20:0] zext_ln50_11_fu_19610_p1;
wire   [20:0] zext_ln50_12_fu_19769_p1;
wire   [20:0] zext_ln50_13_fu_19786_p1;
wire   [20:0] zext_ln50_14_fu_19945_p1;
wire   [20:0] zext_ln50_15_fu_19962_p1;
wire   [20:0] zext_ln50_16_fu_20121_p1;
wire   [20:0] zext_ln50_17_fu_20138_p1;
wire    ap_block_state66_pp0_stage65_iter0;
wire    ap_CS_fsm_state76;
wire    ap_block_state76_pp0_stage75_iter0;
wire  signed [20:0] sext_ln813_fu_1309_p0;
wire  signed [21:0] sext_ln813_36_fu_1313_p1;
wire  signed [21:0] sext_ln813_fu_1309_p1;
wire   [21:0] add_ln1347_fu_1317_p2;
wire  signed [20:0] add_ln813_fu_1331_p1;
wire   [20:0] add_ln813_fu_1331_p2;
wire   [0:0] tmp_fu_1323_p3;
wire   [0:0] tmp_36_fu_1337_p3;
wire   [0:0] xor_ln895_fu_1345_p2;
wire   [0:0] and_ln895_fu_1351_p2;
wire   [0:0] xor_ln302_fu_1357_p2;
wire   [20:0] select_ln346_fu_1363_p3;
wire  signed [20:0] sext_ln813_37_fu_1379_p0;
wire  signed [21:0] sext_ln813_38_fu_1383_p1;
wire  signed [21:0] sext_ln813_37_fu_1379_p1;
wire   [21:0] add_ln1347_1_fu_1387_p2;
wire  signed [20:0] add_ln813_1_fu_1401_p1;
wire   [20:0] add_ln813_1_fu_1401_p2;
wire   [0:0] tmp_37_fu_1393_p3;
wire   [0:0] tmp_38_fu_1407_p3;
wire   [0:0] xor_ln895_18_fu_1415_p2;
wire   [0:0] and_ln895_18_fu_1421_p2;
wire   [0:0] xor_ln302_18_fu_1427_p2;
wire   [20:0] select_ln346_18_fu_1433_p3;
wire  signed [20:0] select_ln302_fu_1371_p3;
wire  signed [20:0] select_ln302_18_fu_1441_p3;
wire  signed [20:0] sext_ln813_39_fu_1457_p0;
wire  signed [21:0] sext_ln813_40_fu_1461_p1;
wire  signed [21:0] sext_ln813_39_fu_1457_p1;
wire   [21:0] add_ln1347_2_fu_1465_p2;
wire  signed [20:0] add_ln813_2_fu_1479_p1;
wire   [20:0] add_ln813_2_fu_1479_p2;
wire   [0:0] tmp_39_fu_1471_p3;
wire   [0:0] tmp_40_fu_1485_p3;
wire   [0:0] xor_ln895_19_fu_1493_p2;
wire   [0:0] and_ln895_19_fu_1499_p2;
wire   [0:0] xor_ln302_19_fu_1505_p2;
wire   [20:0] select_ln346_19_fu_1511_p3;
wire  signed [20:0] sext_ln813_43_fu_1527_p0;
wire  signed [21:0] sext_ln813_44_fu_1531_p1;
wire  signed [21:0] sext_ln813_43_fu_1527_p1;
wire   [21:0] add_ln1347_4_fu_1535_p2;
wire  signed [20:0] add_ln813_4_fu_1549_p1;
wire   [20:0] add_ln813_4_fu_1549_p2;
wire   [0:0] tmp_43_fu_1541_p3;
wire   [0:0] tmp_44_fu_1555_p3;
wire   [0:0] xor_ln895_21_fu_1563_p2;
wire   [0:0] and_ln895_21_fu_1569_p2;
wire   [0:0] xor_ln302_4_fu_1575_p2;
wire   [20:0] select_ln346_21_fu_1581_p3;
wire   [20:0] select_ln302_2_fu_1519_p3;
wire  signed [20:0] select_ln302_19_fu_1589_p3;
wire  signed [20:0] sext_ln813_41_fu_1609_p0;
wire  signed [21:0] sext_ln813_42_fu_1613_p1;
wire  signed [21:0] sext_ln813_41_fu_1609_p1;
wire   [21:0] add_ln1347_3_fu_1617_p2;
wire  signed [20:0] add_ln813_3_fu_1631_p1;
wire   [20:0] add_ln813_3_fu_1631_p2;
wire   [0:0] tmp_41_fu_1623_p3;
wire   [0:0] tmp_42_fu_1637_p3;
wire   [0:0] xor_ln895_20_fu_1645_p2;
wire   [0:0] and_ln895_20_fu_1651_p2;
wire   [0:0] xor_ln302_20_fu_1657_p2;
wire   [20:0] select_ln346_20_fu_1663_p3;
wire  signed [20:0] sext_ln813_45_fu_1679_p0;
wire  signed [21:0] sext_ln813_46_fu_1683_p1;
wire  signed [21:0] sext_ln813_45_fu_1679_p1;
wire   [21:0] add_ln1347_5_fu_1687_p2;
wire  signed [20:0] add_ln813_5_fu_1701_p1;
wire   [20:0] add_ln813_5_fu_1701_p2;
wire   [0:0] tmp_45_fu_1693_p3;
wire   [0:0] tmp_46_fu_1707_p3;
wire   [0:0] xor_ln895_22_fu_1715_p2;
wire   [0:0] and_ln895_22_fu_1721_p2;
wire   [0:0] xor_ln302_5_fu_1727_p2;
wire   [20:0] select_ln346_22_fu_1733_p3;
wire   [6:0] trunc_ln1273_fu_1753_p1;
wire   [8:0] trunc_ln1273_6_fu_1765_p1;
wire   [13:0] trunc_ln1273_1_fu_1769_p3;
wire   [13:0] trunc_ln2_fu_1757_p3;
wire   [13:0] sub_ln1347_fu_1777_p2;
wire   [6:0] trunc_ln1273_7_fu_1799_p1;
wire   [8:0] trunc_ln1273_8_fu_1811_p1;
wire   [13:0] trunc_ln1273_3_fu_1815_p3;
wire   [13:0] trunc_ln1273_2_fu_1803_p3;
wire   [13:0] sub_ln1347_1_fu_1823_p2;
wire  signed [20:0] sext_ln813_47_fu_1837_p0;
wire  signed [21:0] sext_ln813_48_fu_1841_p1;
wire  signed [21:0] sext_ln813_47_fu_1837_p1;
wire   [21:0] add_ln1347_6_fu_1845_p2;
wire  signed [20:0] add_ln813_6_fu_1859_p1;
wire   [20:0] add_ln813_6_fu_1859_p2;
wire   [0:0] tmp_47_fu_1851_p3;
wire   [0:0] tmp_48_fu_1865_p3;
wire   [0:0] xor_ln895_23_fu_1873_p2;
wire   [0:0] and_ln895_23_fu_1879_p2;
wire   [0:0] xor_ln302_6_fu_1885_p2;
wire   [20:0] select_ln346_23_fu_1891_p3;
wire  signed [20:0] sext_ln813_49_fu_1907_p0;
wire  signed [21:0] sext_ln813_50_fu_1911_p1;
wire  signed [21:0] sext_ln813_49_fu_1907_p1;
wire   [21:0] add_ln1347_7_fu_1915_p2;
wire  signed [20:0] add_ln813_7_fu_1929_p1;
wire   [20:0] add_ln813_7_fu_1929_p2;
wire   [0:0] tmp_49_fu_1921_p3;
wire   [0:0] tmp_50_fu_1935_p3;
wire   [0:0] xor_ln895_24_fu_1943_p2;
wire   [0:0] and_ln895_24_fu_1949_p2;
wire   [0:0] xor_ln302_7_fu_1955_p2;
wire   [20:0] select_ln346_24_fu_1961_p3;
wire  signed [34:0] grp_fu_21385_p2;
wire   [0:0] tmp_73_fu_2000_p3;
wire   [20:0] zext_ln377_fu_2007_p1;
wire   [20:0] trunc_ln_fu_1984_p4;
wire   [20:0] add_ln377_fu_2011_p2;
wire   [0:0] tmp_74_fu_2017_p3;
wire   [0:0] tmp_72_fu_1993_p3;
wire   [0:0] xor_ln896_fu_2025_p2;
wire   [0:0] xor_ln888_fu_2044_p2;
wire   [0:0] tmp_75_fu_2037_p3;
wire   [0:0] or_ln888_fu_2050_p2;
wire   [0:0] tmp_76_fu_2062_p3;
wire   [0:0] xor_ln890_fu_2069_p2;
wire   [0:0] or_ln890_fu_2075_p2;
wire   [0:0] and_ln378_fu_2031_p2;
wire   [0:0] xor_ln888_1_fu_2056_p2;
wire   [0:0] xor_ln895_27_fu_2093_p2;
wire   [0:0] tmp_71_fu_1977_p3;
wire   [0:0] or_ln895_fu_2099_p2;
wire   [0:0] xor_ln895_28_fu_2105_p2;
wire   [0:0] and_ln890_fu_2081_p2;
wire   [0:0] xor_ln896_1_fu_2117_p2;
wire   [0:0] and_ln891_fu_2087_p2;
wire   [0:0] or_ln896_fu_2123_p2;
wire   [0:0] xor_ln896_26_fu_2129_p2;
wire   [0:0] and_ln895_35_fu_2111_p2;
wire   [0:0] and_ln896_fu_2135_p2;
wire   [0:0] or_ln346_fu_2141_p2;
wire   [20:0] select_ln346_35_fu_2147_p3;
wire  signed [20:0] select_ln302_20_fu_1899_p3;
wire  signed [20:0] select_ln302_7_fu_1969_p3;
wire  signed [20:0] sext_ln813_51_fu_2178_p0;
wire  signed [21:0] sext_ln813_52_fu_2182_p1;
wire  signed [21:0] sext_ln813_51_fu_2178_p1;
wire   [21:0] add_ln1347_8_fu_2186_p2;
wire  signed [20:0] add_ln813_8_fu_2200_p1;
wire   [20:0] add_ln813_8_fu_2200_p2;
wire   [0:0] tmp_51_fu_2192_p3;
wire   [0:0] tmp_52_fu_2206_p3;
wire   [0:0] xor_ln895_25_fu_2214_p2;
wire   [0:0] and_ln895_25_fu_2220_p2;
wire   [0:0] xor_ln302_8_fu_2226_p2;
wire   [20:0] select_ln346_25_fu_2232_p3;
wire  signed [20:0] sext_ln813_53_fu_2248_p0;
wire  signed [21:0] sext_ln813_54_fu_2252_p1;
wire  signed [21:0] sext_ln813_53_fu_2248_p1;
wire   [21:0] add_ln1347_9_fu_2256_p2;
wire  signed [20:0] add_ln813_9_fu_2270_p1;
wire   [20:0] add_ln813_9_fu_2270_p2;
wire   [0:0] tmp_53_fu_2262_p3;
wire   [0:0] tmp_54_fu_2276_p3;
wire   [0:0] xor_ln895_26_fu_2284_p2;
wire   [0:0] and_ln895_26_fu_2290_p2;
wire   [0:0] xor_ln302_9_fu_2296_p2;
wire   [20:0] select_ln346_26_fu_2302_p3;
wire  signed [34:0] shl_ln_fu_2318_p3;
wire  signed [35:0] sext_ln813_74_fu_2325_p1;
wire  signed [35:0] sext_ln1347_fu_2329_p1;
wire  signed [34:0] sext_ln1347_1_fu_2332_p1;
wire   [35:0] add_ln1347_18_fu_2335_p2;
wire   [34:0] add_ln810_fu_2341_p2;
wire   [20:0] zext_ln377_1_fu_2373_p1;
wire   [20:0] trunc_ln818_1_fu_2355_p4;
wire   [20:0] add_ln377_1_fu_2376_p2;
wire   [0:0] tmp_80_fu_2382_p3;
wire   [0:0] tmp_78_fu_2365_p3;
wire   [0:0] xor_ln896_2_fu_2390_p2;
wire   [0:0] xor_ln888_2_fu_2410_p2;
wire   [0:0] tmp_81_fu_2402_p3;
wire   [0:0] or_ln888_1_fu_2416_p2;
wire   [0:0] tmp_82_fu_2428_p3;
wire   [0:0] xor_ln890_1_fu_2436_p2;
wire   [0:0] or_ln890_1_fu_2442_p2;
wire   [0:0] and_ln378_1_fu_2396_p2;
wire   [0:0] xor_ln888_3_fu_2422_p2;
wire   [0:0] xor_ln895_29_fu_2460_p2;
wire   [0:0] tmp_77_fu_2347_p3;
wire   [0:0] or_ln895_1_fu_2466_p2;
wire   [0:0] xor_ln895_30_fu_2472_p2;
wire   [0:0] and_ln890_1_fu_2448_p2;
wire   [0:0] xor_ln896_3_fu_2484_p2;
wire   [0:0] and_ln891_1_fu_2454_p2;
wire   [0:0] or_ln896_1_fu_2490_p2;
wire   [0:0] xor_ln896_27_fu_2496_p2;
wire   [0:0] and_ln895_36_fu_2478_p2;
wire   [0:0] and_ln896_1_fu_2502_p2;
wire   [0:0] or_ln346_1_fu_2508_p2;
wire   [20:0] select_ln346_37_fu_2514_p3;
wire   [20:0] select_ln302_8_fu_2240_p3;
wire  signed [34:0] grp_fu_21418_p2;
wire   [0:0] tmp_165_fu_2575_p3;
wire   [20:0] zext_ln377_14_fu_2582_p1;
wire   [20:0] trunc_ln818_13_fu_2559_p4;
wire   [20:0] add_ln377_14_fu_2586_p2;
wire   [0:0] tmp_166_fu_2592_p3;
wire   [0:0] tmp_164_fu_2568_p3;
wire   [0:0] xor_ln896_32_fu_2600_p2;
wire   [0:0] xor_ln888_28_fu_2619_p2;
wire   [0:0] tmp_167_fu_2612_p3;
wire   [0:0] or_ln888_14_fu_2625_p2;
wire   [0:0] tmp_168_fu_2637_p3;
wire   [0:0] xor_ln890_14_fu_2644_p2;
wire   [0:0] or_ln890_14_fu_2650_p2;
wire   [0:0] and_ln378_14_fu_2606_p2;
wire   [0:0] xor_ln888_29_fu_2631_p2;
wire   [0:0] xor_ln895_59_fu_2668_p2;
wire   [0:0] tmp_163_fu_2552_p3;
wire   [0:0] or_ln895_14_fu_2674_p2;
wire   [0:0] xor_ln895_60_fu_2680_p2;
wire   [0:0] and_ln890_14_fu_2656_p2;
wire   [0:0] xor_ln896_33_fu_2692_p2;
wire   [0:0] and_ln891_14_fu_2662_p2;
wire   [0:0] or_ln896_14_fu_2698_p2;
wire   [0:0] xor_ln896_70_fu_2704_p2;
wire   [0:0] and_ln895_53_fu_2686_p2;
wire   [0:0] and_ln896_14_fu_2710_p2;
wire   [0:0] or_ln346_14_fu_2716_p2;
wire   [20:0] select_ln346_71_fu_2722_p3;
wire  signed [34:0] grp_fu_21437_p2;
wire   [0:0] tmp_237_fu_2768_p3;
wire   [20:0] zext_ln377_24_fu_2775_p1;
wire   [20:0] trunc_ln818_23_fu_2752_p4;
wire   [20:0] add_ln377_24_fu_2779_p2;
wire   [0:0] tmp_238_fu_2785_p3;
wire   [0:0] tmp_236_fu_2761_p3;
wire   [0:0] xor_ln896_58_fu_2793_p2;
wire   [0:0] xor_ln888_48_fu_2812_p2;
wire   [0:0] tmp_239_fu_2805_p3;
wire   [0:0] or_ln888_24_fu_2818_p2;
wire   [0:0] tmp_240_fu_2830_p3;
wire   [0:0] xor_ln890_24_fu_2837_p2;
wire   [0:0] or_ln890_24_fu_2843_p2;
wire   [0:0] and_ln378_24_fu_2799_p2;
wire   [0:0] xor_ln888_49_fu_2824_p2;
wire   [0:0] xor_ln895_85_fu_2861_p2;
wire   [0:0] tmp_235_fu_2745_p3;
wire   [0:0] or_ln895_24_fu_2867_p2;
wire   [0:0] xor_ln895_86_fu_2873_p2;
wire   [0:0] and_ln890_24_fu_2849_p2;
wire   [0:0] xor_ln896_59_fu_2885_p2;
wire   [0:0] and_ln891_24_fu_2855_p2;
wire   [0:0] or_ln896_24_fu_2891_p2;
wire   [0:0] xor_ln896_128_fu_2897_p2;
wire   [0:0] and_ln895_69_fu_2879_p2;
wire   [0:0] and_ln896_24_fu_2903_p2;
wire   [0:0] or_ln346_24_fu_2909_p2;
wire   [20:0] select_ln346_103_fu_2915_p3;
wire  signed [20:0] sext_ln813_55_fu_2931_p0;
wire  signed [21:0] sext_ln813_56_fu_2935_p1;
wire  signed [21:0] sext_ln813_55_fu_2931_p1;
wire   [21:0] add_ln1347_10_fu_2939_p2;
wire  signed [20:0] add_ln813_10_fu_2953_p1;
wire   [20:0] add_ln813_10_fu_2953_p2;
wire   [0:0] tmp_55_fu_2945_p3;
wire   [0:0] tmp_56_fu_2959_p3;
wire   [0:0] xor_ln895_10_fu_2967_p2;
wire   [0:0] and_ln895_27_fu_2973_p2;
wire   [0:0] xor_ln302_10_fu_2979_p2;
wire   [20:0] select_ln346_27_fu_2985_p3;
wire  signed [20:0] sext_ln813_57_fu_3001_p0;
wire  signed [21:0] sext_ln813_58_fu_3005_p1;
wire  signed [21:0] sext_ln813_57_fu_3001_p1;
wire   [21:0] add_ln1347_11_fu_3009_p2;
wire  signed [20:0] add_ln813_11_fu_3023_p1;
wire   [20:0] add_ln813_11_fu_3023_p2;
wire   [0:0] tmp_57_fu_3015_p3;
wire   [0:0] tmp_58_fu_3029_p3;
wire   [0:0] xor_ln895_11_fu_3037_p2;
wire   [0:0] and_ln895_28_fu_3043_p2;
wire   [0:0] xor_ln302_11_fu_3049_p2;
wire   [20:0] select_ln346_28_fu_3055_p3;
wire  signed [34:0] shl_ln838_1_fu_3071_p3;
wire  signed [35:0] sext_ln813_75_fu_3078_p1;
wire  signed [35:0] sext_ln1347_2_fu_3082_p1;
wire   [35:0] add_ln1347_19_fu_3085_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_1_fu_3091_p2;
wire   [20:0] zext_ln377_2_fu_3122_p1;
wire   [20:0] trunc_ln818_2_fu_3104_p4;
wire   [20:0] add_ln377_2_fu_3125_p2;
wire   [0:0] tmp_86_fu_3131_p3;
wire   [0:0] tmp_84_fu_3114_p3;
wire   [0:0] xor_ln896_4_fu_3139_p2;
wire   [0:0] xor_ln888_4_fu_3159_p2;
wire   [0:0] tmp_87_fu_3151_p3;
wire   [0:0] or_ln888_2_fu_3165_p2;
wire   [0:0] tmp_88_fu_3177_p3;
wire   [0:0] xor_ln890_2_fu_3185_p2;
wire   [0:0] or_ln890_2_fu_3191_p2;
wire   [0:0] and_ln378_2_fu_3145_p2;
wire   [0:0] xor_ln888_5_fu_3171_p2;
wire   [0:0] xor_ln895_31_fu_3209_p2;
wire   [0:0] tmp_83_fu_3096_p3;
wire   [0:0] or_ln895_2_fu_3215_p2;
wire   [0:0] xor_ln895_32_fu_3221_p2;
wire   [0:0] and_ln890_2_fu_3197_p2;
wire   [0:0] xor_ln896_5_fu_3233_p2;
wire   [0:0] and_ln891_2_fu_3203_p2;
wire   [0:0] or_ln896_2_fu_3239_p2;
wire   [0:0] xor_ln896_30_fu_3245_p2;
wire   [0:0] and_ln895_37_fu_3227_p2;
wire   [0:0] and_ln896_2_fu_3251_p2;
wire   [0:0] or_ln346_2_fu_3257_p2;
wire   [20:0] select_ln346_39_fu_3263_p3;
wire  signed [20:0] select_ln302_10_fu_2993_p3;
wire  signed [34:0] shl_ln838_12_fu_3302_p3;
wire  signed [27:0] grp_fu_21456_p2;
wire  signed [35:0] sext_ln813_87_fu_3309_p1;
wire  signed [35:0] sext_ln1347_19_fu_3313_p1;
wire  signed [34:0] sext_ln1347_20_fu_3316_p1;
wire   [35:0] add_ln1347_31_fu_3319_p2;
wire   [34:0] add_ln810_11_fu_3325_p2;
wire   [0:0] tmp_171_fu_3357_p3;
wire   [20:0] zext_ln377_15_fu_3364_p1;
wire   [20:0] trunc_ln818_14_fu_3339_p4;
wire   [0:0] tmp_172_fu_3374_p3;
wire   [0:0] xor_ln888_30_fu_3396_p2;
wire   [0:0] or_ln888_15_fu_3402_p2;
wire   [0:0] tmp_174_fu_3414_p3;
wire   [0:0] xor_ln890_15_fu_3422_p2;
wire   [0:0] or_ln890_15_fu_3428_p2;
wire   [0:0] xor_ln888_31_fu_3408_p2;
wire   [0:0] xor_ln895_61_fu_3440_p2;
wire   [0:0] or_ln895_15_fu_3446_p2;
wire   [0:0] xor_ln895_62_fu_3452_p2;
wire   [0:0] and_ln890_15_fu_3434_p2;
wire   [0:0] xor_ln896_35_fu_3464_p2;
wire  signed [34:0] shl_ln838_21_fu_3476_p3;
wire  signed [27:0] grp_fu_21465_p2;
wire  signed [35:0] sext_ln813_96_fu_3483_p1;
wire  signed [35:0] sext_ln1347_30_fu_3487_p1;
wire  signed [34:0] sext_ln1347_31_fu_3490_p1;
wire   [35:0] add_ln1347_40_fu_3493_p2;
wire   [34:0] add_ln810_18_fu_3499_p2;
wire   [0:0] tmp_243_fu_3531_p3;
wire   [20:0] zext_ln377_25_fu_3538_p1;
wire   [20:0] trunc_ln818_24_fu_3513_p4;
wire   [0:0] tmp_244_fu_3548_p3;
wire   [0:0] xor_ln888_50_fu_3570_p2;
wire   [0:0] or_ln888_25_fu_3576_p2;
wire   [0:0] tmp_246_fu_3588_p3;
wire   [0:0] xor_ln890_25_fu_3596_p2;
wire   [0:0] or_ln890_25_fu_3602_p2;
wire   [0:0] xor_ln888_51_fu_3582_p2;
wire   [0:0] xor_ln895_87_fu_3614_p2;
wire   [0:0] or_ln895_25_fu_3620_p2;
wire   [0:0] xor_ln895_88_fu_3626_p2;
wire   [0:0] and_ln890_25_fu_3608_p2;
wire   [0:0] xor_ln896_61_fu_3638_p2;
wire  signed [20:0] sext_ln813_59_fu_3650_p0;
wire  signed [21:0] sext_ln813_60_fu_3654_p1;
wire  signed [21:0] sext_ln813_59_fu_3650_p1;
wire   [21:0] add_ln1347_12_fu_3658_p2;
wire  signed [20:0] add_ln813_12_fu_3672_p1;
wire   [20:0] add_ln813_12_fu_3672_p2;
wire   [0:0] tmp_59_fu_3664_p3;
wire   [0:0] tmp_60_fu_3678_p3;
wire   [0:0] xor_ln895_12_fu_3686_p2;
wire   [0:0] and_ln895_29_fu_3692_p2;
wire   [0:0] xor_ln302_12_fu_3698_p2;
wire   [20:0] select_ln346_29_fu_3704_p3;
wire  signed [20:0] sext_ln813_61_fu_3720_p0;
wire  signed [21:0] sext_ln813_62_fu_3724_p1;
wire  signed [21:0] sext_ln813_61_fu_3720_p1;
wire   [21:0] add_ln1347_13_fu_3728_p2;
wire  signed [20:0] add_ln813_13_fu_3742_p1;
wire   [20:0] add_ln813_13_fu_3742_p2;
wire   [0:0] tmp_61_fu_3734_p3;
wire   [0:0] tmp_62_fu_3748_p3;
wire   [0:0] xor_ln895_13_fu_3756_p2;
wire   [0:0] and_ln895_30_fu_3762_p2;
wire   [0:0] xor_ln302_13_fu_3768_p2;
wire   [20:0] select_ln346_30_fu_3774_p3;
wire   [27:0] shl_ln1_fu_3790_p3;
wire   [25:0] shl_ln1273_1_fu_3801_p3;
wire  signed [28:0] sext_ln1273_5_fu_3808_p1;
wire  signed [28:0] sext_ln1273_4_fu_3797_p1;
wire  signed [34:0] shl_ln838_2_fu_3818_p3;
wire  signed [28:0] sub_ln1273_fu_3812_p2;
wire  signed [35:0] sext_ln813_76_fu_3825_p1;
wire  signed [35:0] sext_ln1347_3_fu_3829_p1;
wire  signed [34:0] sext_ln1347_4_fu_3833_p1;
wire   [35:0] add_ln1347_20_fu_3837_p2;
wire   [34:0] add_ln810_2_fu_3843_p2;
wire   [20:0] zext_ln377_3_fu_3875_p1;
wire   [20:0] trunc_ln818_3_fu_3857_p4;
wire   [0:0] tmp_92_fu_3884_p3;
wire   [0:0] tmp_90_fu_3867_p3;
wire   [0:0] xor_ln896_6_fu_3892_p2;
wire   [0:0] xor_ln888_6_fu_3912_p2;
wire   [0:0] tmp_93_fu_3904_p3;
wire   [0:0] or_ln888_3_fu_3918_p2;
wire   [0:0] tmp_94_fu_3930_p3;
wire   [0:0] xor_ln890_3_fu_3938_p2;
wire   [0:0] or_ln890_3_fu_3944_p2;
wire   [0:0] and_ln378_3_fu_3898_p2;
wire   [0:0] xor_ln888_7_fu_3924_p2;
wire   [0:0] xor_ln895_33_fu_3962_p2;
wire   [0:0] tmp_89_fu_3849_p3;
wire   [0:0] or_ln895_3_fu_3968_p2;
wire   [0:0] xor_ln895_34_fu_3974_p2;
wire   [0:0] and_ln890_3_fu_3950_p2;
wire   [0:0] xor_ln896_7_fu_3986_p2;
wire   [0:0] and_ln891_3_fu_3956_p2;
wire   [0:0] or_ln896_3_fu_3992_p2;
wire   [0:0] xor_ln896_31_fu_3998_p2;
wire   [0:0] and_ln896_3_fu_4004_p2;
wire  signed [20:0] select_ln302_12_fu_3712_p3;
wire   [0:0] and_ln378_15_fu_4034_p2;
wire   [0:0] and_ln891_15_fu_4038_p2;
wire   [0:0] xor_ln896_71_fu_4043_p2;
wire   [0:0] and_ln896_15_fu_4048_p2;
wire   [0:0] or_ln346_15_fu_4053_p2;
wire   [20:0] select_ln346_73_fu_4058_p3;
wire   [20:0] select_ln346_74_fu_4065_p3;
wire  signed [34:0] shl_ln838_13_fu_4072_p3;
wire  signed [35:0] sext_ln813_88_fu_4080_p1;
wire  signed [35:0] sext_ln1347_21_fu_4084_p1;
wire   [35:0] add_ln1347_32_fu_4087_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_12_fu_4093_p2;
wire   [20:0] zext_ln377_16_fu_4124_p1;
wire   [20:0] trunc_ln818_15_fu_4106_p4;
wire   [0:0] tmp_178_fu_4133_p3;
wire   [0:0] tmp_176_fu_4116_p3;
wire   [0:0] xor_ln896_36_fu_4141_p2;
wire   [0:0] xor_ln888_32_fu_4161_p2;
wire   [0:0] tmp_179_fu_4153_p3;
wire   [0:0] or_ln888_16_fu_4167_p2;
wire   [0:0] tmp_180_fu_4179_p3;
wire   [0:0] xor_ln890_16_fu_4187_p2;
wire   [0:0] or_ln890_16_fu_4193_p2;
wire   [0:0] and_ln378_16_fu_4147_p2;
wire   [0:0] xor_ln888_33_fu_4173_p2;
wire   [0:0] xor_ln895_63_fu_4211_p2;
wire   [0:0] tmp_175_fu_4098_p3;
wire   [0:0] or_ln895_16_fu_4217_p2;
wire   [0:0] xor_ln895_64_fu_4223_p2;
wire   [0:0] and_ln890_16_fu_4199_p2;
wire   [0:0] xor_ln896_37_fu_4235_p2;
wire   [0:0] and_ln891_16_fu_4205_p2;
wire   [0:0] or_ln896_16_fu_4241_p2;
wire   [0:0] xor_ln896_74_fu_4247_p2;
wire   [0:0] and_ln896_16_fu_4253_p2;
wire  signed [20:0] select_ln302_13_fu_3782_p3;
wire   [0:0] and_ln378_25_fu_4269_p2;
wire   [0:0] and_ln891_25_fu_4273_p2;
wire   [0:0] xor_ln896_129_fu_4278_p2;
wire   [0:0] and_ln896_25_fu_4283_p2;
wire   [0:0] or_ln346_25_fu_4295_p2;
wire   [20:0] select_ln346_105_fu_4288_p3;
wire   [20:0] select_ln346_106_fu_4300_p3;
wire   [0:0] tmp_247_fu_4307_p3;
wire   [0:0] tmp_248_fu_4315_p3;
wire   [0:0] xor_ln895_89_fu_4323_p2;
wire   [0:0] and_ln895_71_fu_4329_p2;
wire   [0:0] xor_ln346_10_fu_4343_p2;
wire   [20:0] select_ln346_107_fu_4335_p3;
wire   [20:0] select_ln346_108_fu_4349_p3;
wire   [0:0] tmp_249_fu_4357_p3;
wire   [0:0] tmp_250_fu_4365_p3;
wire   [0:0] xor_ln895_90_fu_4373_p2;
wire   [0:0] and_ln895_72_fu_4379_p2;
wire   [0:0] xor_ln346_11_fu_4393_p2;
wire   [20:0] select_ln346_109_fu_4385_p3;
wire   [20:0] select_ln346_110_fu_4399_p3;
wire   [0:0] tmp_251_fu_4407_p3;
wire   [0:0] tmp_252_fu_4415_p3;
wire   [0:0] xor_ln895_91_fu_4423_p2;
wire   [0:0] and_ln895_73_fu_4429_p2;
wire   [0:0] xor_ln346_12_fu_4443_p2;
wire   [20:0] select_ln346_111_fu_4435_p3;
wire   [20:0] select_ln346_112_fu_4449_p3;
wire   [0:0] tmp_253_fu_4457_p3;
wire   [0:0] tmp_254_fu_4465_p3;
wire   [0:0] xor_ln895_92_fu_4473_p2;
wire   [0:0] and_ln895_74_fu_4479_p2;
wire   [0:0] xor_ln346_13_fu_4485_p2;
wire   [20:0] select_ln346_113_fu_4491_p3;
wire  signed [20:0] sext_ln813_63_fu_4507_p0;
wire  signed [21:0] sext_ln813_64_fu_4511_p1;
wire  signed [21:0] sext_ln813_63_fu_4507_p1;
wire   [21:0] add_ln1347_14_fu_4515_p2;
wire  signed [20:0] add_ln813_14_fu_4529_p1;
wire   [20:0] add_ln813_14_fu_4529_p2;
wire   [0:0] tmp_63_fu_4521_p3;
wire   [0:0] tmp_64_fu_4535_p3;
wire   [0:0] xor_ln895_14_fu_4543_p2;
wire   [0:0] and_ln895_31_fu_4549_p2;
wire   [0:0] xor_ln302_14_fu_4555_p2;
wire   [20:0] select_ln346_31_fu_4561_p3;
wire  signed [20:0] sext_ln813_65_fu_4577_p0;
wire  signed [21:0] sext_ln813_66_fu_4581_p1;
wire  signed [21:0] sext_ln813_65_fu_4577_p1;
wire   [21:0] add_ln1347_15_fu_4585_p2;
wire  signed [20:0] add_ln813_15_fu_4599_p1;
wire   [20:0] add_ln813_15_fu_4599_p2;
wire   [0:0] tmp_65_fu_4591_p3;
wire   [0:0] tmp_66_fu_4605_p3;
wire   [0:0] xor_ln895_15_fu_4613_p2;
wire   [0:0] and_ln895_32_fu_4619_p2;
wire   [0:0] xor_ln302_15_fu_4625_p2;
wire   [20:0] select_ln346_32_fu_4631_p3;
wire   [20:0] select_ln346_41_fu_4647_p3;
wire   [20:0] select_ln346_42_fu_4654_p3;
wire  signed [34:0] shl_ln838_3_fu_4660_p3;
wire  signed [35:0] sext_ln813_77_fu_4668_p1;
wire  signed [35:0] sext_ln1347_5_fu_4672_p1;
wire  signed [34:0] sext_ln1347_6_fu_4675_p1;
wire   [35:0] add_ln1347_21_fu_4678_p2;
wire   [34:0] add_ln810_3_fu_4684_p2;
wire   [20:0] zext_ln377_4_fu_4716_p1;
wire   [20:0] trunc_ln818_4_fu_4698_p4;
wire   [20:0] add_ln377_4_fu_4719_p2;
wire   [0:0] tmp_98_fu_4725_p3;
wire   [0:0] tmp_96_fu_4708_p3;
wire   [0:0] xor_ln896_8_fu_4733_p2;
wire   [0:0] xor_ln888_8_fu_4753_p2;
wire   [0:0] tmp_99_fu_4745_p3;
wire   [0:0] or_ln888_4_fu_4759_p2;
wire   [0:0] tmp_100_fu_4771_p3;
wire   [0:0] xor_ln890_4_fu_4779_p2;
wire   [0:0] or_ln890_4_fu_4785_p2;
wire   [0:0] and_ln378_4_fu_4739_p2;
wire   [0:0] xor_ln888_9_fu_4765_p2;
wire   [0:0] xor_ln895_35_fu_4803_p2;
wire   [0:0] tmp_95_fu_4690_p3;
wire   [0:0] or_ln895_4_fu_4809_p2;
wire   [0:0] xor_ln895_36_fu_4815_p2;
wire   [0:0] and_ln890_4_fu_4791_p2;
wire   [0:0] xor_ln896_9_fu_4827_p2;
wire   [0:0] and_ln891_4_fu_4797_p2;
wire   [0:0] or_ln896_4_fu_4833_p2;
wire   [0:0] xor_ln896_40_fu_4839_p2;
wire   [0:0] and_ln895_39_fu_4821_p2;
wire   [0:0] and_ln896_4_fu_4845_p2;
wire   [0:0] or_ln346_4_fu_4851_p2;
wire   [20:0] select_ln346_43_fu_4857_p3;
wire  signed [20:0] select_ln302_15_fu_4639_p3;
wire   [27:0] shl_ln1273_4_fu_4884_p3;
wire   [25:0] shl_ln1273_5_fu_4895_p3;
wire  signed [28:0] sext_ln1273_23_fu_4902_p1;
wire  signed [28:0] sext_ln1273_22_fu_4891_p1;
wire   [20:0] select_ln346_75_fu_4912_p3;
wire   [20:0] select_ln346_76_fu_4919_p3;
wire  signed [34:0] shl_ln838_14_fu_4925_p3;
wire  signed [28:0] sub_ln1273_2_fu_4906_p2;
wire  signed [35:0] sext_ln813_89_fu_4933_p1;
wire  signed [35:0] sext_ln1347_22_fu_4937_p1;
wire  signed [34:0] sext_ln1347_23_fu_4941_p1;
wire   [35:0] add_ln1347_33_fu_4945_p2;
wire   [34:0] add_ln810_13_fu_4951_p2;
wire   [20:0] zext_ln377_17_fu_4983_p1;
wire   [20:0] trunc_ln818_16_fu_4965_p4;
wire   [0:0] tmp_184_fu_4992_p3;
wire   [0:0] tmp_182_fu_4975_p3;
wire   [0:0] xor_ln896_38_fu_5000_p2;
wire   [0:0] xor_ln888_34_fu_5020_p2;
wire   [0:0] tmp_185_fu_5012_p3;
wire   [0:0] or_ln888_17_fu_5026_p2;
wire   [0:0] tmp_186_fu_5038_p3;
wire   [0:0] xor_ln890_17_fu_5046_p2;
wire   [0:0] or_ln890_17_fu_5052_p2;
wire   [0:0] and_ln378_17_fu_5006_p2;
wire   [0:0] xor_ln888_35_fu_5032_p2;
wire   [0:0] xor_ln895_65_fu_5070_p2;
wire   [0:0] tmp_181_fu_4957_p3;
wire   [0:0] or_ln895_17_fu_5076_p2;
wire   [0:0] xor_ln895_66_fu_5082_p2;
wire   [0:0] and_ln890_17_fu_5058_p2;
wire   [0:0] xor_ln896_39_fu_5094_p2;
wire   [0:0] and_ln891_17_fu_5064_p2;
wire   [0:0] or_ln896_17_fu_5100_p2;
wire   [0:0] xor_ln896_75_fu_5106_p2;
wire   [0:0] and_ln896_17_fu_5112_p2;
wire  signed [20:0] select_ln302_14_fu_4569_p3;
wire  signed [20:0] sext_ln813_67_fu_5142_p0;
wire  signed [21:0] sext_ln813_68_fu_5146_p1;
wire  signed [21:0] sext_ln813_67_fu_5142_p1;
wire   [21:0] add_ln1347_16_fu_5150_p2;
wire  signed [20:0] add_ln813_16_fu_5164_p1;
wire   [20:0] add_ln813_16_fu_5164_p2;
wire   [0:0] tmp_67_fu_5156_p3;
wire   [0:0] tmp_68_fu_5170_p3;
wire   [0:0] xor_ln895_16_fu_5178_p2;
wire   [0:0] and_ln895_33_fu_5184_p2;
wire   [0:0] xor_ln302_16_fu_5190_p2;
wire   [20:0] select_ln346_33_fu_5196_p3;
wire  signed [20:0] sext_ln813_69_fu_5212_p0;
wire  signed [21:0] sext_ln813_70_fu_5216_p1;
wire  signed [21:0] sext_ln813_69_fu_5212_p1;
wire   [21:0] add_ln1347_17_fu_5220_p2;
wire  signed [20:0] add_ln813_17_fu_5234_p1;
wire   [20:0] add_ln813_17_fu_5234_p2;
wire   [0:0] tmp_69_fu_5226_p3;
wire   [0:0] tmp_70_fu_5240_p3;
wire   [0:0] xor_ln895_17_fu_5248_p2;
wire   [0:0] and_ln895_34_fu_5254_p2;
wire   [0:0] xor_ln302_17_fu_5260_p2;
wire   [20:0] select_ln346_34_fu_5266_p3;
wire  signed [34:0] shl_ln838_4_fu_5282_p3;
wire  signed [35:0] sext_ln813_78_fu_5289_p1;
wire  signed [35:0] sext_ln1347_7_fu_5293_p1;
wire  signed [34:0] sext_ln1347_8_fu_5296_p1;
wire   [35:0] add_ln1347_22_fu_5299_p2;
wire   [34:0] add_ln810_4_fu_5305_p2;
wire   [20:0] zext_ln377_5_fu_5337_p1;
wire   [20:0] trunc_ln818_5_fu_5319_p4;
wire   [20:0] add_ln377_5_fu_5340_p2;
wire   [0:0] tmp_104_fu_5346_p3;
wire   [0:0] tmp_102_fu_5329_p3;
wire   [0:0] xor_ln896_10_fu_5354_p2;
wire   [0:0] xor_ln888_10_fu_5374_p2;
wire   [0:0] tmp_105_fu_5366_p3;
wire   [0:0] or_ln888_5_fu_5380_p2;
wire   [0:0] tmp_106_fu_5392_p3;
wire   [0:0] xor_ln890_5_fu_5400_p2;
wire   [0:0] or_ln890_5_fu_5406_p2;
wire   [0:0] and_ln378_5_fu_5360_p2;
wire   [0:0] xor_ln888_11_fu_5386_p2;
wire   [0:0] xor_ln895_37_fu_5424_p2;
wire   [0:0] tmp_101_fu_5311_p3;
wire   [0:0] or_ln895_5_fu_5430_p2;
wire   [0:0] xor_ln895_38_fu_5436_p2;
wire   [0:0] and_ln890_5_fu_5412_p2;
wire   [0:0] xor_ln896_11_fu_5448_p2;
wire   [0:0] and_ln891_5_fu_5418_p2;
wire   [0:0] or_ln896_5_fu_5454_p2;
wire   [0:0] xor_ln896_41_fu_5460_p2;
wire   [0:0] and_ln895_40_fu_5442_p2;
wire   [0:0] and_ln896_5_fu_5466_p2;
wire   [0:0] or_ln346_5_fu_5472_p2;
wire   [20:0] select_ln346_45_fu_5478_p3;
wire   [20:0] select_ln346_77_fu_5508_p3;
wire   [20:0] select_ln346_78_fu_5515_p3;
wire   [0:0] tmp_187_fu_5521_p3;
wire   [0:0] tmp_188_fu_5529_p3;
wire   [0:0] xor_ln895_67_fu_5537_p2;
wire   [0:0] and_ln895_57_fu_5543_p2;
wire   [0:0] xor_ln346_4_fu_5557_p2;
wire   [20:0] select_ln346_79_fu_5549_p3;
wire   [20:0] select_ln346_80_fu_5563_p3;
wire   [0:0] tmp_189_fu_5571_p3;
wire   [0:0] tmp_190_fu_5579_p3;
wire   [0:0] xor_ln895_68_fu_5587_p2;
wire   [0:0] and_ln895_58_fu_5593_p2;
wire   [0:0] xor_ln346_5_fu_5599_p2;
wire   [20:0] select_ln346_81_fu_5605_p3;
wire   [20:0] select_ln346_82_fu_5613_p3;
wire  signed [34:0] shl_ln838_15_fu_5621_p3;
wire  signed [35:0] sext_ln813_90_fu_5629_p1;
wire  signed [35:0] sext_ln1347_24_fu_5633_p1;
wire   [35:0] add_ln1347_34_fu_5636_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_14_fu_5642_p2;
wire   [20:0] zext_ln377_18_fu_5673_p1;
wire   [20:0] trunc_ln818_17_fu_5655_p4;
wire   [0:0] tmp_194_fu_5682_p3;
wire   [0:0] xor_ln888_36_fu_5704_p2;
wire   [0:0] or_ln888_18_fu_5710_p2;
wire   [0:0] tmp_196_fu_5722_p3;
wire   [0:0] xor_ln890_18_fu_5730_p2;
wire   [0:0] or_ln890_18_fu_5736_p2;
wire   [0:0] xor_ln888_37_fu_5716_p2;
wire   [0:0] xor_ln895_69_fu_5748_p2;
wire   [0:0] or_ln895_18_fu_5754_p2;
wire   [0:0] xor_ln895_70_fu_5760_p2;
wire   [0:0] and_ln890_18_fu_5742_p2;
wire   [0:0] xor_ln896_43_fu_5772_p2;
wire  signed [20:0] select_ln302_16_fu_5204_p3;
wire  signed [34:0] shl_ln838_22_fu_5795_p3;
wire  signed [34:0] grp_fu_21530_p2;
wire  signed [35:0] sext_ln813_97_fu_5802_p1;
wire  signed [35:0] sext_ln1347_32_fu_5806_p1;
wire   [35:0] add_ln1347_41_fu_5809_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_19_fu_5815_p2;
wire   [0:0] tmp_257_fu_5846_p3;
wire   [20:0] zext_ln377_26_fu_5853_p1;
wire   [20:0] trunc_ln818_25_fu_5828_p4;
wire   [0:0] tmp_258_fu_5863_p3;
wire   [0:0] xor_ln888_52_fu_5885_p2;
wire   [0:0] or_ln888_26_fu_5891_p2;
wire   [0:0] tmp_260_fu_5903_p3;
wire   [0:0] xor_ln890_26_fu_5911_p2;
wire   [0:0] or_ln890_26_fu_5917_p2;
wire   [0:0] xor_ln888_53_fu_5897_p2;
wire   [0:0] xor_ln895_93_fu_5929_p2;
wire   [0:0] or_ln895_26_fu_5935_p2;
wire   [0:0] xor_ln895_94_fu_5941_p2;
wire   [0:0] and_ln890_26_fu_5923_p2;
wire   [0:0] xor_ln896_67_fu_5953_p2;
wire  signed [20:0] select_ln302_17_fu_5274_p3;
wire  signed [34:0] shl_ln838_5_fu_5976_p3;
wire  signed [35:0] sext_ln813_79_fu_5983_p1;
wire  signed [35:0] sext_ln1347_9_fu_5987_p1;
wire   [35:0] add_ln1347_23_fu_5990_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_5_fu_5996_p2;
wire   [20:0] zext_ln377_6_fu_6027_p1;
wire   [20:0] trunc_ln818_6_fu_6009_p4;
wire   [20:0] add_ln377_6_fu_6030_p2;
wire   [0:0] tmp_110_fu_6036_p3;
wire   [0:0] tmp_108_fu_6019_p3;
wire   [0:0] xor_ln896_12_fu_6044_p2;
wire   [0:0] xor_ln888_12_fu_6064_p2;
wire   [0:0] tmp_111_fu_6056_p3;
wire   [0:0] or_ln888_6_fu_6070_p2;
wire   [0:0] tmp_112_fu_6082_p3;
wire   [0:0] xor_ln890_6_fu_6090_p2;
wire   [0:0] or_ln890_6_fu_6096_p2;
wire   [0:0] and_ln378_6_fu_6050_p2;
wire   [0:0] xor_ln888_13_fu_6076_p2;
wire   [0:0] xor_ln895_39_fu_6114_p2;
wire   [0:0] tmp_107_fu_6001_p3;
wire   [0:0] or_ln895_6_fu_6120_p2;
wire   [0:0] xor_ln895_40_fu_6126_p2;
wire   [0:0] and_ln890_6_fu_6102_p2;
wire   [0:0] xor_ln896_13_fu_6138_p2;
wire   [0:0] and_ln891_6_fu_6108_p2;
wire   [0:0] or_ln896_6_fu_6144_p2;
wire   [0:0] xor_ln896_50_fu_6150_p2;
wire   [0:0] and_ln895_41_fu_6132_p2;
wire   [0:0] and_ln896_6_fu_6156_p2;
wire   [0:0] or_ln346_6_fu_6162_p2;
wire   [20:0] select_ln346_47_fu_6168_p3;
wire   [0:0] and_ln378_18_fu_6191_p2;
wire   [0:0] and_ln891_18_fu_6195_p2;
wire   [0:0] xor_ln896_98_fu_6200_p2;
wire   [0:0] and_ln896_18_fu_6205_p2;
wire   [0:0] or_ln346_18_fu_6210_p2;
wire   [20:0] select_ln346_83_fu_6215_p3;
wire   [20:0] select_ln346_84_fu_6222_p3;
wire  signed [34:0] shl_ln838_16_fu_6229_p3;
wire  signed [35:0] sext_ln813_91_fu_6237_p1;
wire  signed [35:0] sext_ln1347_25_fu_6241_p1;
wire  signed [34:0] sext_ln1347_26_fu_6244_p1;
wire   [35:0] add_ln1347_35_fu_6247_p2;
wire   [34:0] add_ln810_15_fu_6253_p2;
wire   [20:0] zext_ln377_19_fu_6285_p1;
wire   [20:0] trunc_ln818_18_fu_6267_p4;
wire   [0:0] tmp_200_fu_6294_p3;
wire   [0:0] tmp_198_fu_6277_p3;
wire   [0:0] xor_ln896_44_fu_6302_p2;
wire   [0:0] xor_ln888_38_fu_6322_p2;
wire   [0:0] tmp_201_fu_6314_p3;
wire   [0:0] or_ln888_19_fu_6328_p2;
wire   [0:0] tmp_202_fu_6340_p3;
wire   [0:0] xor_ln890_19_fu_6348_p2;
wire   [0:0] or_ln890_19_fu_6354_p2;
wire   [0:0] and_ln378_19_fu_6308_p2;
wire   [0:0] xor_ln888_39_fu_6334_p2;
wire   [0:0] xor_ln895_71_fu_6372_p2;
wire   [0:0] tmp_197_fu_6259_p3;
wire   [0:0] or_ln895_19_fu_6378_p2;
wire   [0:0] xor_ln895_72_fu_6384_p2;
wire   [0:0] and_ln890_19_fu_6360_p2;
wire   [0:0] xor_ln896_45_fu_6396_p2;
wire   [0:0] and_ln891_19_fu_6366_p2;
wire   [0:0] or_ln896_19_fu_6402_p2;
wire   [0:0] xor_ln896_99_fu_6408_p2;
wire   [0:0] and_ln896_19_fu_6414_p2;
wire   [0:0] and_ln378_26_fu_6433_p2;
wire   [0:0] and_ln891_26_fu_6437_p2;
wire   [0:0] xor_ln896_132_fu_6442_p2;
wire   [0:0] and_ln896_26_fu_6447_p2;
wire   [0:0] or_ln346_26_fu_6452_p2;
wire   [20:0] select_ln346_115_fu_6457_p3;
wire   [20:0] select_ln346_116_fu_6464_p3;
wire  signed [34:0] shl_ln838_23_fu_6471_p3;
wire  signed [35:0] sext_ln813_98_fu_6479_p1;
wire  signed [35:0] sext_ln1347_33_fu_6483_p1;
wire  signed [34:0] sext_ln1347_34_fu_6486_p1;
wire   [35:0] add_ln1347_42_fu_6489_p2;
wire   [34:0] add_ln810_20_fu_6495_p2;
wire   [20:0] zext_ln377_27_fu_6527_p1;
wire   [20:0] trunc_ln818_26_fu_6509_p4;
wire   [0:0] tmp_264_fu_6536_p3;
wire   [0:0] tmp_262_fu_6519_p3;
wire   [0:0] xor_ln896_68_fu_6544_p2;
wire   [0:0] xor_ln888_54_fu_6564_p2;
wire   [0:0] tmp_265_fu_6556_p3;
wire   [0:0] or_ln888_27_fu_6570_p2;
wire   [0:0] tmp_266_fu_6582_p3;
wire   [0:0] xor_ln890_27_fu_6590_p2;
wire   [0:0] or_ln890_27_fu_6596_p2;
wire   [0:0] and_ln378_27_fu_6550_p2;
wire   [0:0] xor_ln888_55_fu_6576_p2;
wire   [0:0] xor_ln895_95_fu_6614_p2;
wire   [0:0] tmp_261_fu_6501_p3;
wire   [0:0] or_ln895_27_fu_6620_p2;
wire   [0:0] xor_ln895_96_fu_6626_p2;
wire   [0:0] and_ln890_27_fu_6602_p2;
wire   [0:0] xor_ln896_69_fu_6638_p2;
wire   [0:0] and_ln891_27_fu_6608_p2;
wire   [0:0] or_ln896_27_fu_6644_p2;
wire   [0:0] xor_ln896_133_fu_6650_p2;
wire   [0:0] and_ln896_27_fu_6656_p2;
wire  signed [34:0] shl_ln838_6_fu_6668_p3;
wire  signed [35:0] sext_ln813_80_fu_6675_p1;
wire  signed [35:0] sext_ln1347_10_fu_6679_p1;
wire  signed [34:0] sext_ln1347_11_fu_6682_p1;
wire   [35:0] add_ln1347_24_fu_6685_p2;
wire   [34:0] add_ln810_6_fu_6691_p2;
wire   [20:0] zext_ln377_7_fu_6723_p1;
wire   [20:0] trunc_ln818_7_fu_6705_p4;
wire   [20:0] add_ln377_7_fu_6726_p2;
wire   [0:0] tmp_116_fu_6732_p3;
wire   [0:0] tmp_114_fu_6715_p3;
wire   [0:0] xor_ln896_14_fu_6740_p2;
wire   [0:0] xor_ln888_14_fu_6760_p2;
wire   [0:0] tmp_117_fu_6752_p3;
wire   [0:0] or_ln888_7_fu_6766_p2;
wire   [0:0] tmp_118_fu_6778_p3;
wire   [0:0] xor_ln890_7_fu_6786_p2;
wire   [0:0] or_ln890_7_fu_6792_p2;
wire   [0:0] and_ln378_7_fu_6746_p2;
wire   [0:0] xor_ln888_15_fu_6772_p2;
wire   [0:0] xor_ln895_41_fu_6810_p2;
wire   [0:0] tmp_113_fu_6697_p3;
wire   [0:0] or_ln895_7_fu_6816_p2;
wire   [0:0] xor_ln895_42_fu_6822_p2;
wire   [0:0] and_ln890_7_fu_6798_p2;
wire   [0:0] xor_ln896_15_fu_6834_p2;
wire   [0:0] and_ln891_7_fu_6804_p2;
wire   [0:0] or_ln896_7_fu_6840_p2;
wire   [0:0] xor_ln896_53_fu_6846_p2;
wire   [0:0] and_ln895_42_fu_6828_p2;
wire   [0:0] and_ln896_7_fu_6852_p2;
wire   [0:0] or_ln346_7_fu_6858_p2;
wire   [20:0] select_ln346_49_fu_6864_p3;
wire   [20:0] select_ln346_85_fu_6887_p3;
wire   [20:0] select_ln346_86_fu_6894_p3;
wire  signed [34:0] shl_ln838_17_fu_6900_p3;
wire  signed [35:0] sext_ln813_92_fu_6908_p1;
wire  signed [35:0] sext_ln1347_27_fu_6912_p1;
wire   [35:0] add_ln1347_36_fu_6915_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_16_fu_6921_p2;
wire   [20:0] zext_ln377_20_fu_6952_p1;
wire   [20:0] trunc_ln818_19_fu_6934_p4;
wire   [20:0] add_ln377_20_fu_6955_p2;
wire   [0:0] tmp_206_fu_6961_p3;
wire   [0:0] tmp_204_fu_6944_p3;
wire   [0:0] xor_ln896_46_fu_6969_p2;
wire   [0:0] xor_ln888_40_fu_6989_p2;
wire   [0:0] tmp_207_fu_6981_p3;
wire   [0:0] or_ln888_20_fu_6995_p2;
wire   [0:0] tmp_208_fu_7007_p3;
wire   [0:0] xor_ln890_20_fu_7015_p2;
wire   [0:0] or_ln890_20_fu_7021_p2;
wire   [0:0] and_ln378_20_fu_6975_p2;
wire   [0:0] xor_ln888_41_fu_7001_p2;
wire   [0:0] xor_ln895_73_fu_7039_p2;
wire   [0:0] tmp_203_fu_6926_p3;
wire   [0:0] or_ln895_20_fu_7045_p2;
wire   [0:0] xor_ln895_74_fu_7051_p2;
wire   [0:0] and_ln890_20_fu_7027_p2;
wire   [0:0] xor_ln896_47_fu_7063_p2;
wire   [0:0] and_ln891_20_fu_7033_p2;
wire   [0:0] or_ln896_20_fu_7069_p2;
wire   [0:0] xor_ln896_102_fu_7075_p2;
wire   [0:0] and_ln895_61_fu_7057_p2;
wire   [0:0] and_ln896_20_fu_7081_p2;
wire   [0:0] or_ln346_20_fu_7087_p2;
wire   [20:0] select_ln346_87_fu_7093_p3;
wire   [20:0] select_ln346_117_fu_7109_p3;
wire   [20:0] select_ln346_118_fu_7116_p3;
wire   [0:0] tmp_267_fu_7122_p3;
wire   [0:0] tmp_268_fu_7130_p3;
wire   [0:0] xor_ln895_97_fu_7138_p2;
wire   [0:0] and_ln895_77_fu_7144_p2;
wire   [0:0] xor_ln346_14_fu_7158_p2;
wire   [20:0] select_ln346_119_fu_7150_p3;
wire   [20:0] select_ln346_120_fu_7164_p3;
wire   [0:0] tmp_269_fu_7172_p3;
wire   [0:0] tmp_270_fu_7180_p3;
wire   [0:0] xor_ln895_98_fu_7188_p2;
wire   [0:0] and_ln895_78_fu_7194_p2;
wire   [0:0] xor_ln346_15_fu_7200_p2;
wire   [20:0] select_ln346_121_fu_7206_p3;
wire   [20:0] select_ln346_122_fu_7214_p3;
wire   [34:0] shl_ln838_24_fu_7222_p3;
wire  signed [35:0] sext_ln813_99_fu_7230_p1;
wire  signed [35:0] grp_fu_21567_p2;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_43_fu_7234_p2;
wire   [0:0] tmp_273_fu_7265_p3;
wire   [20:0] zext_ln377_28_fu_7272_p1;
wire   [20:0] trunc_ln818_27_fu_7247_p4;
wire   [0:0] tmp_274_fu_7282_p3;
wire   [0:0] xor_ln888_56_fu_7304_p2;
wire   [0:0] or_ln888_28_fu_7310_p2;
wire   [0:0] tmp_276_fu_7322_p3;
wire   [0:0] xor_ln890_28_fu_7330_p2;
wire   [0:0] or_ln890_28_fu_7336_p2;
wire   [0:0] xor_ln888_57_fu_7316_p2;
wire   [0:0] xor_ln895_99_fu_7348_p2;
wire   [0:0] or_ln895_28_fu_7354_p2;
wire   [0:0] xor_ln895_100_fu_7360_p2;
wire   [0:0] and_ln890_28_fu_7342_p2;
wire   [0:0] xor_ln896_73_fu_7372_p2;
wire  signed [34:0] shl_ln838_7_fu_7384_p3;
wire  signed [35:0] sext_ln813_81_fu_7391_p1;
wire  signed [35:0] sext_ln1347_12_fu_7395_p1;
wire   [35:0] add_ln1347_25_fu_7398_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_7_fu_7404_p2;
wire   [20:0] zext_ln377_8_fu_7435_p1;
wire   [20:0] trunc_ln818_8_fu_7417_p4;
wire   [20:0] add_ln377_8_fu_7438_p2;
wire   [0:0] tmp_122_fu_7444_p3;
wire   [0:0] tmp_120_fu_7427_p3;
wire   [0:0] xor_ln896_16_fu_7452_p2;
wire   [0:0] xor_ln888_16_fu_7472_p2;
wire   [0:0] tmp_123_fu_7464_p3;
wire   [0:0] or_ln888_8_fu_7478_p2;
wire   [0:0] tmp_124_fu_7490_p3;
wire   [0:0] xor_ln890_8_fu_7498_p2;
wire   [0:0] or_ln890_8_fu_7504_p2;
wire   [0:0] and_ln378_8_fu_7458_p2;
wire   [0:0] xor_ln888_17_fu_7484_p2;
wire   [0:0] xor_ln895_43_fu_7522_p2;
wire   [0:0] tmp_119_fu_7409_p3;
wire   [0:0] or_ln895_8_fu_7528_p2;
wire   [0:0] xor_ln895_44_fu_7534_p2;
wire   [0:0] and_ln890_8_fu_7510_p2;
wire   [0:0] xor_ln896_17_fu_7546_p2;
wire   [0:0] and_ln891_8_fu_7516_p2;
wire   [0:0] or_ln896_8_fu_7552_p2;
wire   [0:0] xor_ln896_54_fu_7558_p2;
wire   [0:0] and_ln895_43_fu_7540_p2;
wire   [0:0] and_ln896_8_fu_7564_p2;
wire   [0:0] or_ln346_8_fu_7570_p2;
wire   [20:0] select_ln346_51_fu_7576_p3;
wire   [27:0] shl_ln1273_6_fu_7592_p3;
wire   [25:0] shl_ln1273_7_fu_7603_p3;
wire  signed [28:0] sext_ln1273_24_fu_7599_p1;
wire  signed [28:0] sext_ln1273_25_fu_7610_p1;
wire  signed [34:0] shl_ln838_18_fu_7620_p3;
wire  signed [28:0] sub_ln1273_3_fu_7614_p2;
wire  signed [35:0] sext_ln813_93_fu_7627_p1;
wire  signed [35:0] sext_ln1347_28_fu_7631_p1;
wire  signed [34:0] sext_ln1347_29_fu_7635_p1;
wire   [35:0] add_ln1347_37_fu_7639_p2;
wire   [34:0] add_ln810_17_fu_7645_p2;
wire   [0:0] tmp_211_fu_7677_p3;
wire   [20:0] zext_ln377_21_fu_7685_p1;
wire   [20:0] trunc_ln818_20_fu_7659_p4;
wire   [0:0] tmp_212_fu_7695_p3;
wire   [0:0] tmp_210_fu_7669_p3;
wire   [0:0] xor_ln896_48_fu_7703_p2;
wire   [0:0] xor_ln888_42_fu_7723_p2;
wire   [0:0] tmp_213_fu_7715_p3;
wire   [0:0] or_ln888_21_fu_7729_p2;
wire   [0:0] tmp_214_fu_7741_p3;
wire   [0:0] xor_ln890_21_fu_7749_p2;
wire   [0:0] or_ln890_21_fu_7755_p2;
wire   [0:0] and_ln378_21_fu_7709_p2;
wire   [0:0] xor_ln888_43_fu_7735_p2;
wire   [0:0] xor_ln895_75_fu_7773_p2;
wire   [0:0] tmp_209_fu_7651_p3;
wire   [0:0] or_ln895_21_fu_7779_p2;
wire   [0:0] xor_ln895_76_fu_7785_p2;
wire   [0:0] and_ln890_21_fu_7761_p2;
wire   [0:0] xor_ln896_49_fu_7797_p2;
wire   [0:0] and_ln891_21_fu_7767_p2;
wire   [0:0] or_ln896_21_fu_7803_p2;
wire   [0:0] xor_ln896_103_fu_7809_p2;
wire   [0:0] and_ln896_21_fu_7815_p2;
wire   [0:0] and_ln378_28_fu_7834_p2;
wire   [0:0] and_ln891_28_fu_7838_p2;
wire   [0:0] xor_ln896_138_fu_7843_p2;
wire   [0:0] and_ln896_28_fu_7848_p2;
wire   [0:0] or_ln346_28_fu_7860_p2;
wire   [20:0] select_ln346_123_fu_7853_p3;
wire   [20:0] select_ln346_124_fu_7865_p3;
wire   [0:0] tmp_277_fu_7872_p3;
wire   [0:0] tmp_278_fu_7880_p3;
wire   [0:0] xor_ln895_101_fu_7888_p2;
wire   [0:0] and_ln895_80_fu_7894_p2;
wire   [0:0] xor_ln346_16_fu_7908_p2;
wire   [20:0] select_ln346_125_fu_7900_p3;
wire   [20:0] select_ln346_126_fu_7914_p3;
wire   [0:0] tmp_279_fu_7922_p3;
wire   [0:0] tmp_280_fu_7930_p3;
wire   [0:0] xor_ln895_102_fu_7938_p2;
wire   [0:0] and_ln895_81_fu_7944_p2;
wire   [0:0] xor_ln346_17_fu_7950_p2;
wire   [20:0] select_ln346_127_fu_7956_p3;
wire   [20:0] select_ln346_128_fu_7964_p3;
wire   [34:0] shl_ln838_25_fu_7972_p3;
wire  signed [35:0] sext_ln813_101_fu_7980_p1;
wire  signed [35:0] grp_fu_21582_p2;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_44_fu_7984_p2;
wire   [0:0] tmp_283_fu_8015_p3;
wire   [20:0] zext_ln377_29_fu_8022_p1;
wire   [20:0] trunc_ln818_28_fu_7997_p4;
wire   [0:0] tmp_284_fu_8032_p3;
wire   [0:0] xor_ln888_58_fu_8054_p2;
wire   [0:0] or_ln888_29_fu_8060_p2;
wire   [0:0] tmp_286_fu_8072_p3;
wire   [0:0] xor_ln890_29_fu_8080_p2;
wire   [0:0] or_ln890_29_fu_8086_p2;
wire   [0:0] xor_ln888_59_fu_8066_p2;
wire   [0:0] xor_ln895_103_fu_8098_p2;
wire   [0:0] or_ln895_29_fu_8104_p2;
wire   [0:0] xor_ln895_104_fu_8110_p2;
wire   [0:0] and_ln890_29_fu_8092_p2;
wire   [0:0] xor_ln896_77_fu_8122_p2;
wire   [27:0] shl_ln1273_2_fu_8134_p3;
wire   [25:0] shl_ln1273_3_fu_8145_p3;
wire  signed [28:0] sext_ln1273_14_fu_8141_p1;
wire  signed [28:0] sext_ln1273_15_fu_8152_p1;
wire  signed [34:0] shl_ln838_8_fu_8162_p3;
wire  signed [28:0] sub_ln1273_1_fu_8156_p2;
wire  signed [35:0] sext_ln813_82_fu_8169_p1;
wire  signed [35:0] sext_ln1347_13_fu_8173_p1;
wire  signed [34:0] sext_ln1347_14_fu_8177_p1;
wire   [35:0] add_ln1347_26_fu_8181_p2;
wire   [34:0] add_ln810_8_fu_8187_p2;
wire   [0:0] tmp_127_fu_8219_p3;
wire   [20:0] zext_ln377_9_fu_8227_p1;
wire   [20:0] trunc_ln818_9_fu_8201_p4;
wire   [0:0] tmp_128_fu_8237_p3;
wire   [0:0] tmp_126_fu_8211_p3;
wire   [0:0] xor_ln896_18_fu_8245_p2;
wire   [0:0] xor_ln888_18_fu_8265_p2;
wire   [0:0] tmp_129_fu_8257_p3;
wire   [0:0] or_ln888_9_fu_8271_p2;
wire   [0:0] tmp_130_fu_8283_p3;
wire   [0:0] xor_ln890_9_fu_8291_p2;
wire   [0:0] or_ln890_9_fu_8297_p2;
wire   [0:0] and_ln378_9_fu_8251_p2;
wire   [0:0] xor_ln888_19_fu_8277_p2;
wire   [0:0] xor_ln895_45_fu_8315_p2;
wire   [0:0] tmp_125_fu_8193_p3;
wire   [0:0] or_ln895_9_fu_8321_p2;
wire   [0:0] xor_ln895_46_fu_8327_p2;
wire   [0:0] and_ln890_9_fu_8303_p2;
wire   [0:0] xor_ln896_19_fu_8339_p2;
wire   [0:0] and_ln891_9_fu_8309_p2;
wire   [0:0] or_ln896_9_fu_8345_p2;
wire   [0:0] xor_ln896_57_fu_8351_p2;
wire   [0:0] and_ln896_9_fu_8357_p2;
wire   [20:0] select_ln346_89_fu_8369_p3;
wire   [20:0] select_ln346_90_fu_8376_p3;
wire   [0:0] tmp_215_fu_8382_p3;
wire   [0:0] tmp_216_fu_8390_p3;
wire   [0:0] xor_ln895_77_fu_8398_p2;
wire   [0:0] and_ln895_63_fu_8404_p2;
wire   [0:0] xor_ln346_6_fu_8410_p2;
wire   [20:0] select_ln346_91_fu_8416_p3;
wire   [20:0] select_ln346_92_fu_8424_p3;
wire   [34:0] shl_ln838_19_fu_8432_p3;
wire  signed [35:0] sext_ln813_94_fu_8440_p1;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_38_fu_8444_p2;
wire   [20:0] zext_ln377_22_fu_8475_p1;
wire   [20:0] trunc_ln818_21_fu_8457_p4;
wire   [0:0] tmp_220_fu_8484_p3;
wire   [0:0] tmp_218_fu_8467_p3;
wire   [0:0] xor_ln896_51_fu_8492_p2;
wire   [0:0] xor_ln888_44_fu_8512_p2;
wire   [0:0] tmp_221_fu_8504_p3;
wire   [0:0] or_ln888_22_fu_8518_p2;
wire   [0:0] tmp_222_fu_8530_p3;
wire   [0:0] xor_ln890_22_fu_8538_p2;
wire   [0:0] or_ln890_22_fu_8544_p2;
wire   [0:0] and_ln378_22_fu_8498_p2;
wire   [0:0] xor_ln888_45_fu_8524_p2;
wire   [0:0] xor_ln895_78_fu_8562_p2;
wire   [0:0] tmp_217_fu_8449_p3;
wire   [0:0] or_ln895_22_fu_8568_p2;
wire   [0:0] xor_ln895_79_fu_8574_p2;
wire   [0:0] and_ln890_22_fu_8550_p2;
wire   [0:0] xor_ln896_52_fu_8586_p2;
wire   [0:0] and_ln891_22_fu_8556_p2;
wire   [0:0] or_ln896_22_fu_8592_p2;
wire   [0:0] xor_ln896_108_fu_8598_p2;
wire   [0:0] and_ln896_22_fu_8604_p2;
wire   [0:0] and_ln378_29_fu_8616_p2;
wire   [0:0] and_ln891_29_fu_8620_p2;
wire   [0:0] xor_ln896_143_fu_8625_p2;
wire   [0:0] and_ln896_29_fu_8630_p2;
wire   [0:0] or_ln346_29_fu_8642_p2;
wire   [20:0] select_ln346_129_fu_8635_p3;
wire   [20:0] select_ln346_130_fu_8647_p3;
wire  signed [21:0] sext_ln813_103_fu_8654_p1;
wire   [21:0] sub_ln1348_19_fu_8658_p2;
wire   [0:0] tmp_291_fu_8663_p3;
wire   [0:0] tmp_292_fu_8675_p3;
wire   [0:0] xor_ln895_107_fu_8683_p2;
wire   [0:0] and_ln895_85_fu_8689_p2;
wire   [0:0] xor_ln302_23_fu_8695_p2;
wire   [20:0] select_ln346_133_fu_8701_p3;
wire   [20:0] trunc_ln813_19_fu_8671_p1;
wire  signed [20:0] select_ln302_23_fu_8709_p3;
wire   [28:0] shl_ln1273_8_fu_8725_p3;
wire   [5:0] trunc_ln1273_9_fu_8737_p1;
wire  signed [29:0] sext_ln1273_38_fu_8733_p1;
wire   [13:0] trunc_ln1273_10_fu_8749_p1;
wire   [13:0] trunc_ln1273_4_fu_8741_p3;
wire   [13:0] sub_ln1347_2_fu_8759_p2;
wire   [20:0] select_ln346_53_fu_8773_p3;
wire   [20:0] select_ln346_54_fu_8780_p3;
wire  signed [34:0] shl_ln838_9_fu_8786_p3;
wire  signed [35:0] sext_ln813_83_fu_8794_p1;
wire  signed [35:0] sext_ln1347_15_fu_8798_p1;
wire  signed [34:0] sext_ln1347_16_fu_8801_p1;
wire   [35:0] add_ln1347_27_fu_8804_p2;
wire   [34:0] add_ln810_9_fu_8810_p2;
wire   [20:0] zext_ln377_10_fu_8842_p1;
wire   [20:0] trunc_ln818_s_fu_8824_p4;
wire   [20:0] add_ln377_10_fu_8845_p2;
wire   [0:0] tmp_134_fu_8851_p3;
wire   [0:0] tmp_132_fu_8834_p3;
wire   [0:0] xor_ln896_20_fu_8859_p2;
wire   [0:0] xor_ln888_20_fu_8879_p2;
wire   [0:0] tmp_135_fu_8871_p3;
wire   [0:0] or_ln888_10_fu_8885_p2;
wire   [0:0] tmp_136_fu_8897_p3;
wire   [0:0] xor_ln890_10_fu_8905_p2;
wire   [0:0] or_ln890_10_fu_8911_p2;
wire   [0:0] and_ln378_10_fu_8865_p2;
wire   [0:0] xor_ln888_21_fu_8891_p2;
wire   [0:0] xor_ln895_47_fu_8929_p2;
wire   [0:0] tmp_131_fu_8816_p3;
wire   [0:0] or_ln895_10_fu_8935_p2;
wire   [0:0] xor_ln895_48_fu_8941_p2;
wire   [0:0] and_ln890_10_fu_8917_p2;
wire   [0:0] xor_ln896_21_fu_8953_p2;
wire   [0:0] and_ln891_10_fu_8923_p2;
wire   [0:0] or_ln896_10_fu_8959_p2;
wire   [0:0] xor_ln896_62_fu_8965_p2;
wire   [0:0] and_ln895_45_fu_8947_p2;
wire   [0:0] and_ln896_10_fu_8971_p2;
wire   [0:0] or_ln346_10_fu_8977_p2;
wire   [20:0] select_ln346_55_fu_8983_p3;
wire   [20:0] select_ln346_93_fu_8999_p3;
wire   [20:0] select_ln346_94_fu_9006_p3;
wire   [0:0] tmp_223_fu_9012_p3;
wire   [0:0] tmp_224_fu_9020_p3;
wire   [0:0] xor_ln895_80_fu_9028_p2;
wire   [0:0] and_ln895_65_fu_9034_p2;
wire   [0:0] xor_ln346_7_fu_9048_p2;
wire   [20:0] select_ln346_95_fu_9040_p3;
wire   [20:0] select_ln346_96_fu_9054_p3;
wire   [0:0] tmp_225_fu_9062_p3;
wire   [0:0] tmp_226_fu_9070_p3;
wire   [0:0] xor_ln895_81_fu_9078_p2;
wire   [0:0] and_ln895_66_fu_9084_p2;
wire   [0:0] xor_ln346_8_fu_9090_p2;
wire   [20:0] select_ln346_97_fu_9096_p3;
wire   [20:0] select_ln346_98_fu_9104_p3;
wire   [34:0] shl_ln838_20_fu_9112_p3;
wire  signed [35:0] sext_ln813_95_fu_9120_p1;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_39_fu_9124_p2;
wire   [20:0] zext_ln377_23_fu_9155_p1;
wire   [20:0] trunc_ln818_22_fu_9137_p4;
wire   [0:0] tmp_230_fu_9164_p3;
wire   [0:0] tmp_228_fu_9147_p3;
wire   [0:0] xor_ln896_55_fu_9172_p2;
wire   [0:0] xor_ln888_46_fu_9192_p2;
wire   [0:0] tmp_231_fu_9184_p3;
wire   [0:0] or_ln888_23_fu_9198_p2;
wire   [0:0] tmp_232_fu_9210_p3;
wire   [0:0] xor_ln890_23_fu_9218_p2;
wire   [0:0] or_ln890_23_fu_9224_p2;
wire   [0:0] and_ln378_23_fu_9178_p2;
wire   [0:0] xor_ln888_47_fu_9204_p2;
wire   [0:0] xor_ln895_82_fu_9242_p2;
wire   [0:0] tmp_227_fu_9129_p3;
wire   [0:0] or_ln895_23_fu_9248_p2;
wire   [0:0] xor_ln895_83_fu_9254_p2;
wire   [0:0] and_ln890_23_fu_9230_p2;
wire   [0:0] xor_ln896_56_fu_9266_p2;
wire   [0:0] and_ln891_23_fu_9236_p2;
wire   [0:0] or_ln896_23_fu_9272_p2;
wire   [0:0] xor_ln896_113_fu_9278_p2;
wire   [0:0] and_ln896_23_fu_9284_p2;
wire  signed [34:0] shl_ln838_s_fu_9296_p3;
wire  signed [35:0] sext_ln813_84_fu_9303_p1;
wire  signed [35:0] sext_ln1347_17_fu_9307_p1;
wire  signed [34:0] sext_ln1347_18_fu_9310_p1;
wire   [35:0] add_ln1347_28_fu_9313_p2;
wire   [34:0] add_ln810_10_fu_9319_p2;
wire   [20:0] zext_ln377_11_fu_9351_p1;
wire   [20:0] trunc_ln818_10_fu_9333_p4;
wire   [0:0] tmp_140_fu_9360_p3;
wire   [0:0] tmp_138_fu_9343_p3;
wire   [0:0] xor_ln896_22_fu_9368_p2;
wire   [0:0] xor_ln888_22_fu_9388_p2;
wire   [0:0] tmp_141_fu_9380_p3;
wire   [0:0] or_ln888_11_fu_9394_p2;
wire   [0:0] tmp_142_fu_9406_p3;
wire   [0:0] xor_ln890_11_fu_9414_p2;
wire   [0:0] or_ln890_11_fu_9420_p2;
wire   [0:0] and_ln378_11_fu_9374_p2;
wire   [0:0] xor_ln888_23_fu_9400_p2;
wire   [0:0] xor_ln895_49_fu_9438_p2;
wire   [0:0] tmp_137_fu_9325_p3;
wire   [0:0] or_ln895_11_fu_9444_p2;
wire   [0:0] xor_ln895_50_fu_9450_p2;
wire   [0:0] and_ln890_11_fu_9426_p2;
wire   [0:0] xor_ln896_23_fu_9462_p2;
wire   [0:0] and_ln891_11_fu_9432_p2;
wire   [0:0] or_ln896_11_fu_9468_p2;
wire   [0:0] xor_ln896_63_fu_9474_p2;
wire   [0:0] and_ln896_11_fu_9480_p2;
wire   [20:0] select_ln346_99_fu_9492_p3;
wire   [20:0] select_ln346_100_fu_9499_p3;
wire   [0:0] tmp_233_fu_9505_p3;
wire   [0:0] tmp_234_fu_9513_p3;
wire   [0:0] xor_ln895_84_fu_9521_p2;
wire   [0:0] and_ln895_68_fu_9527_p2;
wire   [0:0] xor_ln346_9_fu_9541_p2;
wire   [20:0] select_ln346_101_fu_9533_p3;
wire   [20:0] select_ln346_102_fu_9547_p3;
wire  signed [21:0] sext_ln813_102_fu_9555_p1;
wire   [21:0] sub_ln1348_18_fu_9559_p2;
wire   [0:0] tmp_289_fu_9564_p3;
wire   [0:0] tmp_290_fu_9576_p3;
wire   [0:0] xor_ln895_106_fu_9584_p2;
wire   [0:0] and_ln895_84_fu_9590_p2;
wire   [0:0] xor_ln302_22_fu_9596_p2;
wire   [20:0] select_ln346_132_fu_9602_p3;
wire   [20:0] trunc_ln813_18_fu_9572_p1;
wire   [5:0] trunc_ln1273_11_fu_9626_p1;
wire   [13:0] trunc_ln1273_12_fu_9638_p1;
wire   [13:0] trunc_ln1273_5_fu_9630_p3;
wire   [13:0] sub_ln1347_3_fu_9642_p2;
wire   [20:0] select_ln346_57_fu_9656_p3;
wire   [20:0] select_ln346_58_fu_9663_p3;
wire   [34:0] shl_ln838_10_fu_9669_p3;
wire  signed [35:0] sext_ln813_85_fu_9677_p1;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_29_fu_9681_p2;
wire   [20:0] zext_ln377_12_fu_9712_p1;
wire   [20:0] trunc_ln818_11_fu_9694_p4;
wire   [0:0] tmp_146_fu_9721_p3;
wire   [0:0] tmp_144_fu_9704_p3;
wire   [0:0] xor_ln896_24_fu_9729_p2;
wire   [0:0] xor_ln888_24_fu_9749_p2;
wire   [0:0] tmp_147_fu_9741_p3;
wire   [0:0] or_ln888_12_fu_9755_p2;
wire   [0:0] tmp_148_fu_9767_p3;
wire   [0:0] xor_ln890_12_fu_9775_p2;
wire   [0:0] or_ln890_12_fu_9781_p2;
wire   [0:0] and_ln378_12_fu_9735_p2;
wire   [0:0] xor_ln888_25_fu_9761_p2;
wire   [0:0] xor_ln895_51_fu_9799_p2;
wire   [0:0] tmp_143_fu_9686_p3;
wire   [0:0] or_ln895_12_fu_9805_p2;
wire   [0:0] xor_ln895_52_fu_9811_p2;
wire   [0:0] and_ln890_12_fu_9787_p2;
wire   [0:0] xor_ln896_25_fu_9823_p2;
wire   [0:0] and_ln891_12_fu_9793_p2;
wire   [0:0] or_ln896_12_fu_9829_p2;
wire   [0:0] xor_ln896_64_fu_9835_p2;
wire   [0:0] and_ln896_12_fu_9841_p2;
wire   [20:0] select_ln346_59_fu_9867_p3;
wire   [20:0] select_ln346_60_fu_9874_p3;
wire   [0:0] tmp_149_fu_9880_p3;
wire   [0:0] tmp_150_fu_9888_p3;
wire   [0:0] xor_ln895_53_fu_9896_p2;
wire   [0:0] and_ln895_48_fu_9902_p2;
wire   [0:0] xor_ln346_fu_9916_p2;
wire   [20:0] select_ln346_61_fu_9908_p3;
wire   [20:0] select_ln346_62_fu_9922_p3;
wire   [0:0] tmp_151_fu_9930_p3;
wire   [0:0] tmp_152_fu_9938_p3;
wire   [0:0] xor_ln895_54_fu_9946_p2;
wire   [0:0] and_ln895_49_fu_9952_p2;
wire   [0:0] xor_ln346_1_fu_9958_p2;
wire   [20:0] select_ln346_63_fu_9964_p3;
wire   [20:0] select_ln346_64_fu_9972_p3;
wire   [34:0] shl_ln838_11_fu_9980_p3;
wire  signed [35:0] sext_ln813_86_fu_9988_p1;
(* use_dsp48 = "no" *) wire   [35:0] add_ln1347_30_fu_9992_p2;
wire   [20:0] zext_ln377_13_fu_10023_p1;
wire   [20:0] trunc_ln818_12_fu_10005_p4;
wire   [0:0] tmp_156_fu_10032_p3;
wire   [0:0] tmp_154_fu_10015_p3;
wire   [0:0] xor_ln896_28_fu_10040_p2;
wire   [0:0] xor_ln888_26_fu_10060_p2;
wire   [0:0] tmp_157_fu_10052_p3;
wire   [0:0] or_ln888_13_fu_10066_p2;
wire   [0:0] tmp_158_fu_10078_p3;
wire   [0:0] xor_ln890_13_fu_10086_p2;
wire   [0:0] or_ln890_13_fu_10092_p2;
wire   [0:0] and_ln378_13_fu_10046_p2;
wire   [0:0] xor_ln888_27_fu_10072_p2;
wire   [0:0] xor_ln895_55_fu_10110_p2;
wire   [0:0] tmp_153_fu_9997_p3;
wire   [0:0] or_ln895_13_fu_10116_p2;
wire   [0:0] xor_ln895_56_fu_10122_p2;
wire   [0:0] and_ln890_13_fu_10098_p2;
wire   [0:0] xor_ln896_29_fu_10134_p2;
wire   [0:0] and_ln891_13_fu_10104_p2;
wire   [0:0] or_ln896_13_fu_10140_p2;
wire   [0:0] xor_ln896_65_fu_10146_p2;
wire   [0:0] and_ln896_13_fu_10152_p2;
wire   [20:0] select_ln346_65_fu_10164_p3;
wire   [20:0] select_ln346_66_fu_10171_p3;
wire   [0:0] tmp_159_fu_10177_p3;
wire   [0:0] tmp_160_fu_10185_p3;
wire   [0:0] xor_ln895_57_fu_10193_p2;
wire   [0:0] and_ln895_51_fu_10199_p2;
wire   [0:0] xor_ln346_2_fu_10213_p2;
wire   [20:0] select_ln346_67_fu_10205_p3;
wire   [20:0] select_ln346_68_fu_10219_p3;
wire   [0:0] tmp_161_fu_10227_p3;
wire   [0:0] tmp_162_fu_10235_p3;
wire   [0:0] xor_ln895_58_fu_10243_p2;
wire   [0:0] and_ln895_52_fu_10249_p2;
wire   [0:0] xor_ln346_3_fu_10263_p2;
wire   [20:0] select_ln346_69_fu_10255_p3;
wire   [20:0] select_ln346_70_fu_10269_p3;
wire  signed [21:0] sext_ln813_100_fu_10277_p1;
wire   [21:0] sub_ln1348_fu_10281_p2;
wire   [0:0] tmp_287_fu_10286_p3;
wire   [0:0] tmp_288_fu_10298_p3;
wire   [0:0] xor_ln895_105_fu_10306_p2;
wire   [0:0] and_ln895_83_fu_10312_p2;
wire   [0:0] xor_ln302_21_fu_10318_p2;
wire   [20:0] select_ln346_131_fu_10324_p3;
wire   [20:0] trunc_ln813_fu_10294_p1;
wire  signed [20:0] select_ln302_21_fu_10332_p3;
wire  signed [33:0] grp_fu_21618_p2;
wire   [19:0] trunc_ln818_29_fu_10373_p4;
wire   [0:0] tmp_295_fu_10393_p3;
wire   [20:0] zext_ln377_30_fu_10400_p1;
wire  signed [20:0] sext_ln818_fu_10382_p1;
wire   [20:0] add_ln377_30_fu_10404_p2;
wire   [0:0] tmp_296_fu_10410_p3;
wire   [0:0] tmp_294_fu_10386_p3;
wire   [0:0] xor_ln896_78_fu_10418_p2;
wire   [0:0] xor_ln888_60_fu_10437_p2;
wire   [0:0] tmp_297_fu_10430_p3;
wire   [0:0] or_ln888_30_fu_10443_p2;
wire   [0:0] tmp_298_fu_10455_p3;
wire   [0:0] xor_ln890_30_fu_10462_p2;
wire   [0:0] or_ln890_30_fu_10468_p2;
wire   [0:0] and_ln378_30_fu_10424_p2;
wire   [0:0] xor_ln888_61_fu_10449_p2;
wire   [0:0] xor_ln895_108_fu_10486_p2;
wire   [0:0] tmp_293_fu_10366_p3;
wire   [0:0] or_ln895_30_fu_10492_p2;
wire   [0:0] xor_ln895_109_fu_10498_p2;
wire   [0:0] and_ln890_30_fu_10474_p2;
wire   [0:0] xor_ln896_79_fu_10510_p2;
wire   [0:0] and_ln891_30_fu_10480_p2;
wire   [0:0] or_ln896_30_fu_10516_p2;
wire   [0:0] xor_ln896_156_fu_10522_p2;
wire   [0:0] and_ln895_86_fu_10504_p2;
wire   [0:0] and_ln896_30_fu_10528_p2;
wire   [0:0] or_ln346_30_fu_10534_p2;
wire   [20:0] select_ln346_134_fu_10540_p3;
wire  signed [30:0] grp_fu_21630_p2;
wire   [16:0] trunc_ln818_32_fu_10563_p4;
wire   [0:0] tmp_313_fu_10583_p3;
wire   [17:0] zext_ln377_33_fu_10590_p1;
wire  signed [17:0] sext_ln365_fu_10572_p1;
wire   [0:0] tmp_314_fu_10600_p3;
wire   [0:0] tmp_312_fu_10576_p3;
wire   [0:0] xor_ln896_84_fu_10608_p2;
wire   [0:0] xor_ln888_66_fu_10627_p2;
wire   [0:0] tmp_315_fu_10620_p3;
wire   [0:0] or_ln888_33_fu_10633_p2;
wire   [0:0] tmp_316_fu_10645_p3;
wire   [0:0] xor_ln890_33_fu_10652_p2;
wire   [0:0] or_ln890_33_fu_10658_p2;
wire   [0:0] and_ln378_33_fu_10614_p2;
wire   [0:0] xor_ln888_67_fu_10639_p2;
wire   [0:0] xor_ln895_114_fu_10676_p2;
wire   [0:0] tmp_311_fu_10556_p3;
wire   [0:0] or_ln895_33_fu_10682_p2;
wire   [0:0] xor_ln895_115_fu_10688_p2;
wire   [0:0] and_ln890_33_fu_10664_p2;
wire   [0:0] xor_ln896_85_fu_10700_p2;
wire   [0:0] and_ln891_33_fu_10670_p2;
wire   [0:0] or_ln896_33_fu_10706_p2;
wire   [0:0] xor_ln896_160_fu_10712_p2;
wire   [0:0] and_ln896_33_fu_10718_p2;
wire  signed [29:0] grp_fu_21642_p2;
wire   [15:0] trunc_ln818_35_fu_10737_p4;
wire   [0:0] tmp_331_fu_10757_p3;
wire   [16:0] zext_ln377_36_fu_10764_p1;
wire  signed [16:0] sext_ln365_1_fu_10746_p1;
wire   [0:0] tmp_332_fu_10774_p3;
wire   [0:0] tmp_330_fu_10750_p3;
wire   [0:0] xor_ln896_90_fu_10782_p2;
wire   [0:0] xor_ln888_72_fu_10801_p2;
wire   [0:0] tmp_333_fu_10794_p3;
wire   [0:0] or_ln888_36_fu_10807_p2;
wire   [0:0] tmp_334_fu_10819_p3;
wire   [0:0] xor_ln890_36_fu_10826_p2;
wire   [0:0] or_ln890_36_fu_10832_p2;
wire   [0:0] and_ln378_36_fu_10788_p2;
wire   [0:0] xor_ln888_73_fu_10813_p2;
wire   [0:0] xor_ln895_120_fu_10850_p2;
wire   [0:0] tmp_329_fu_10730_p3;
wire   [0:0] or_ln895_36_fu_10856_p2;
wire   [0:0] xor_ln895_121_fu_10862_p2;
wire   [0:0] and_ln890_36_fu_10838_p2;
wire   [0:0] xor_ln896_91_fu_10874_p2;
wire   [0:0] and_ln891_36_fu_10844_p2;
wire   [0:0] or_ln896_36_fu_10880_p2;
wire   [0:0] xor_ln896_164_fu_10886_p2;
wire   [0:0] and_ln896_36_fu_10892_p2;
wire  signed [34:0] shl_ln838_26_fu_10907_p3;
wire  signed [35:0] sext_ln813_104_fu_10914_p1;
wire  signed [35:0] sext_ln1347_35_fu_10918_p1;
wire  signed [34:0] sext_ln1347_36_fu_10921_p1;
wire   [35:0] add_ln1347_45_fu_10924_p2;
wire   [34:0] add_ln810_21_fu_10930_p2;
wire   [20:0] zext_ln377_31_fu_10962_p1;
wire   [20:0] trunc_ln818_30_fu_10944_p4;
wire   [20:0] add_ln377_31_fu_10965_p2;
wire   [0:0] tmp_302_fu_10971_p3;
wire   [0:0] tmp_300_fu_10954_p3;
wire   [0:0] xor_ln896_80_fu_10979_p2;
wire   [0:0] xor_ln888_62_fu_10999_p2;
wire   [0:0] tmp_303_fu_10991_p3;
wire   [0:0] or_ln888_31_fu_11005_p2;
wire   [0:0] tmp_304_fu_11017_p3;
wire   [0:0] xor_ln890_31_fu_11025_p2;
wire   [0:0] or_ln890_31_fu_11031_p2;
wire   [0:0] and_ln378_31_fu_10985_p2;
wire   [0:0] xor_ln888_63_fu_11011_p2;
wire   [0:0] xor_ln895_110_fu_11049_p2;
wire   [0:0] tmp_299_fu_10936_p3;
wire   [0:0] or_ln895_31_fu_11055_p2;
wire   [0:0] xor_ln895_111_fu_11061_p2;
wire   [0:0] and_ln890_31_fu_11037_p2;
wire   [0:0] xor_ln896_81_fu_11073_p2;
wire   [0:0] and_ln891_31_fu_11043_p2;
wire   [0:0] or_ln896_31_fu_11079_p2;
wire   [0:0] xor_ln896_157_fu_11085_p2;
wire   [0:0] and_ln895_87_fu_11067_p2;
wire   [0:0] and_ln896_31_fu_11091_p2;
wire   [0:0] or_ln346_31_fu_11097_p2;
wire   [20:0] select_ln346_136_fu_11103_p3;
wire   [20:0] select_ln346_140_fu_11122_p3;
wire  signed [20:0] sext_ln856_fu_11119_p1;
wire   [20:0] select_ln346_141_fu_11129_p3;
wire  signed [34:0] shl_ln838_28_fu_11136_p3;
wire  signed [35:0] sext_ln813_106_fu_11144_p1;
wire  signed [35:0] sext_ln1347_39_fu_11148_p1;
wire  signed [34:0] sext_ln1347_40_fu_11151_p1;
wire   [35:0] add_ln1347_47_fu_11154_p2;
wire   [34:0] add_ln810_23_fu_11160_p2;
wire   [20:0] zext_ln377_34_fu_11192_p1;
wire   [20:0] trunc_ln818_33_fu_11174_p4;
wire   [20:0] add_ln377_34_fu_11195_p2;
wire   [0:0] tmp_320_fu_11201_p3;
wire   [0:0] tmp_318_fu_11184_p3;
wire   [0:0] xor_ln896_86_fu_11209_p2;
wire   [0:0] xor_ln888_68_fu_11229_p2;
wire   [0:0] tmp_321_fu_11221_p3;
wire   [0:0] or_ln888_34_fu_11235_p2;
wire   [0:0] tmp_322_fu_11247_p3;
wire   [0:0] xor_ln890_34_fu_11255_p2;
wire   [0:0] or_ln890_34_fu_11261_p2;
wire   [0:0] and_ln378_34_fu_11215_p2;
wire   [0:0] xor_ln888_69_fu_11241_p2;
wire   [0:0] xor_ln895_116_fu_11279_p2;
wire   [0:0] tmp_317_fu_11166_p3;
wire   [0:0] or_ln895_34_fu_11285_p2;
wire   [0:0] xor_ln895_117_fu_11291_p2;
wire   [0:0] and_ln890_34_fu_11267_p2;
wire   [0:0] xor_ln896_87_fu_11303_p2;
wire   [0:0] and_ln891_34_fu_11273_p2;
wire   [0:0] or_ln896_34_fu_11309_p2;
wire   [0:0] xor_ln896_162_fu_11315_p2;
wire   [0:0] and_ln895_90_fu_11297_p2;
wire   [0:0] and_ln896_34_fu_11321_p2;
wire   [0:0] or_ln346_34_fu_11327_p2;
wire   [20:0] select_ln346_142_fu_11333_p3;
wire   [28:0] shl_ln1273_9_fu_11352_p3;
wire  signed [29:0] sext_ln1273_33_fu_10904_p1;
wire  signed [29:0] sext_ln1273_39_fu_11359_p1;
wire   [20:0] select_ln346_146_fu_11369_p3;
wire  signed [20:0] sext_ln856_1_fu_11349_p1;
wire   [20:0] select_ln346_147_fu_11376_p3;
wire  signed [34:0] shl_ln838_30_fu_11383_p3;
wire  signed [29:0] sub_ln1273_5_fu_11363_p2;
wire  signed [35:0] sext_ln813_108_fu_11391_p1;
wire  signed [35:0] sext_ln1347_43_fu_11395_p1;
wire  signed [34:0] sext_ln1347_44_fu_11399_p1;
wire   [35:0] add_ln1347_49_fu_11403_p2;
wire   [34:0] add_ln810_25_fu_11409_p2;
wire   [20:0] zext_ln377_37_fu_11441_p1;
wire   [20:0] trunc_ln818_36_fu_11423_p4;
wire   [0:0] tmp_338_fu_11450_p3;
wire   [0:0] tmp_336_fu_11433_p3;
wire   [0:0] xor_ln896_92_fu_11458_p2;
wire   [0:0] xor_ln888_74_fu_11478_p2;
wire   [0:0] tmp_339_fu_11470_p3;
wire   [0:0] or_ln888_37_fu_11484_p2;
wire   [0:0] tmp_340_fu_11496_p3;
wire   [0:0] xor_ln890_37_fu_11504_p2;
wire   [0:0] or_ln890_37_fu_11510_p2;
wire   [0:0] and_ln378_37_fu_11464_p2;
wire   [0:0] xor_ln888_75_fu_11490_p2;
wire   [0:0] xor_ln895_122_fu_11528_p2;
wire   [0:0] tmp_335_fu_11415_p3;
wire   [0:0] or_ln895_37_fu_11534_p2;
wire   [0:0] xor_ln895_123_fu_11540_p2;
wire   [0:0] and_ln890_37_fu_11516_p2;
wire   [0:0] xor_ln896_93_fu_11552_p2;
wire   [0:0] and_ln891_37_fu_11522_p2;
wire   [0:0] or_ln896_37_fu_11558_p2;
wire   [0:0] xor_ln896_165_fu_11564_p2;
wire   [0:0] and_ln896_37_fu_11570_p2;
wire  signed [34:0] shl_ln838_27_fu_11582_p3;
wire  signed [35:0] sext_ln813_105_fu_11589_p1;
wire  signed [35:0] sext_ln1347_37_fu_11593_p1;
wire  signed [34:0] sext_ln1347_38_fu_11596_p1;
wire   [35:0] add_ln1347_46_fu_11599_p2;
wire   [34:0] add_ln810_22_fu_11605_p2;
wire   [20:0] zext_ln377_32_fu_11637_p1;
wire   [20:0] trunc_ln818_31_fu_11619_p4;
wire   [0:0] tmp_308_fu_11646_p3;
wire   [0:0] tmp_306_fu_11629_p3;
wire   [0:0] xor_ln896_82_fu_11654_p2;
wire   [0:0] xor_ln888_64_fu_11674_p2;
wire   [0:0] tmp_309_fu_11666_p3;
wire   [0:0] or_ln888_32_fu_11680_p2;
wire   [0:0] tmp_310_fu_11692_p3;
wire   [0:0] xor_ln890_32_fu_11700_p2;
wire   [0:0] or_ln890_32_fu_11706_p2;
wire   [0:0] and_ln378_32_fu_11660_p2;
wire   [0:0] xor_ln888_65_fu_11686_p2;
wire   [0:0] xor_ln895_112_fu_11724_p2;
wire   [0:0] tmp_305_fu_11611_p3;
wire   [0:0] or_ln895_32_fu_11730_p2;
wire   [0:0] xor_ln895_113_fu_11736_p2;
wire   [0:0] and_ln890_32_fu_11712_p2;
wire   [0:0] xor_ln896_83_fu_11748_p2;
wire   [0:0] and_ln891_32_fu_11718_p2;
wire   [0:0] or_ln896_32_fu_11754_p2;
wire   [0:0] xor_ln896_158_fu_11760_p2;
wire   [0:0] and_ln896_32_fu_11766_p2;
wire  signed [34:0] shl_ln838_29_fu_11778_p3;
wire  signed [35:0] sext_ln813_107_fu_11785_p1;
wire  signed [35:0] sext_ln1347_41_fu_11789_p1;
wire  signed [34:0] sext_ln1347_42_fu_11792_p1;
wire   [35:0] add_ln1347_48_fu_11795_p2;
wire   [34:0] add_ln810_24_fu_11801_p2;
wire   [20:0] zext_ln377_35_fu_11833_p1;
wire   [20:0] trunc_ln818_34_fu_11815_p4;
wire   [0:0] tmp_326_fu_11842_p3;
wire   [0:0] tmp_324_fu_11825_p3;
wire   [0:0] xor_ln896_88_fu_11850_p2;
wire   [0:0] xor_ln888_70_fu_11870_p2;
wire   [0:0] tmp_327_fu_11862_p3;
wire   [0:0] or_ln888_35_fu_11876_p2;
wire   [0:0] tmp_328_fu_11888_p3;
wire   [0:0] xor_ln890_35_fu_11896_p2;
wire   [0:0] or_ln890_35_fu_11902_p2;
wire   [0:0] and_ln378_35_fu_11856_p2;
wire   [0:0] xor_ln888_71_fu_11882_p2;
wire   [0:0] xor_ln895_118_fu_11920_p2;
wire   [0:0] tmp_323_fu_11807_p3;
wire   [0:0] or_ln895_35_fu_11926_p2;
wire   [0:0] xor_ln895_119_fu_11932_p2;
wire   [0:0] and_ln890_35_fu_11908_p2;
wire   [0:0] xor_ln896_89_fu_11944_p2;
wire   [0:0] and_ln891_35_fu_11914_p2;
wire   [0:0] or_ln896_35_fu_11950_p2;
wire   [0:0] xor_ln896_163_fu_11956_p2;
wire   [0:0] and_ln896_35_fu_11962_p2;
wire   [20:0] select_ln346_148_fu_11974_p3;
wire   [20:0] select_ln346_149_fu_11981_p3;
wire  signed [34:0] shl_ln838_31_fu_11987_p3;
wire  signed [35:0] sext_ln813_109_fu_11995_p1;
wire  signed [35:0] sext_ln1347_45_fu_11999_p1;
wire   [35:0] add_ln1347_50_fu_12002_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_26_fu_12008_p2;
wire   [20:0] zext_ln377_38_fu_12039_p1;
wire   [20:0] trunc_ln818_37_fu_12021_p4;
wire   [0:0] tmp_344_fu_12048_p3;
wire   [0:0] tmp_342_fu_12031_p3;
wire   [0:0] xor_ln896_94_fu_12056_p2;
wire   [0:0] xor_ln888_76_fu_12076_p2;
wire   [0:0] tmp_345_fu_12068_p3;
wire   [0:0] or_ln888_38_fu_12082_p2;
wire   [0:0] tmp_346_fu_12094_p3;
wire   [0:0] xor_ln890_38_fu_12102_p2;
wire   [0:0] or_ln890_38_fu_12108_p2;
wire   [0:0] and_ln378_38_fu_12062_p2;
wire   [0:0] xor_ln888_77_fu_12088_p2;
wire   [0:0] xor_ln895_124_fu_12126_p2;
wire   [0:0] tmp_341_fu_12013_p3;
wire   [0:0] or_ln895_38_fu_12132_p2;
wire   [0:0] xor_ln895_125_fu_12138_p2;
wire   [0:0] and_ln890_38_fu_12114_p2;
wire   [0:0] xor_ln896_95_fu_12150_p2;
wire   [0:0] and_ln891_38_fu_12120_p2;
wire   [0:0] or_ln896_38_fu_12156_p2;
wire   [0:0] xor_ln896_166_fu_12162_p2;
wire   [0:0] and_ln896_38_fu_12168_p2;
wire   [20:0] select_ln346_138_fu_12180_p3;
wire   [20:0] select_ln346_144_fu_12199_p3;
wire   [0:0] tmp_515_fu_12240_p3;
wire   [0:0] tmp_516_fu_12248_p3;
wire   [0:0] xor_ln895_186_fu_12256_p2;
wire   [0:0] and_ln895_131_fu_12262_p2;
wire   [0:0] xor_ln346_30_fu_12276_p2;
wire   [20:0] select_ln346_224_fu_12268_p3;
wire   [20:0] select_ln346_225_fu_12282_p3;
wire   [0:0] tmp_517_fu_12290_p3;
wire   [0:0] tmp_518_fu_12298_p3;
wire   [0:0] xor_ln895_187_fu_12306_p2;
wire   [0:0] and_ln895_132_fu_12312_p2;
wire   [0:0] xor_ln346_31_fu_12326_p2;
wire   [20:0] select_ln346_226_fu_12318_p3;
wire   [20:0] select_ln346_227_fu_12332_p3;
wire   [0:0] tmp_519_fu_12340_p3;
wire   [0:0] tmp_520_fu_12348_p3;
wire   [0:0] xor_ln895_188_fu_12356_p2;
wire   [0:0] and_ln895_133_fu_12362_p2;
wire   [0:0] xor_ln346_32_fu_12376_p2;
wire   [20:0] select_ln346_228_fu_12368_p3;
wire   [0:0] tmp_522_fu_12399_p3;
wire   [0:0] tmp_523_fu_12407_p3;
wire   [0:0] tmp_521_fu_12391_p3;
wire   [0:0] or_ln895_63_fu_12415_p2;
wire   [0:0] xor_ln895_189_fu_12421_p2;
wire   [0:0] and_ln896_63_fu_12433_p2;
wire   [0:0] xor_ln896_159_fu_12439_p2;
wire   [0:0] and_ln895_134_fu_12427_p2;
wire   [0:0] and_ln896_64_fu_12445_p2;
wire   [0:0] or_ln346_63_fu_12459_p2;
wire   [20:0] select_ln346_230_fu_12451_p3;
wire   [20:0] select_ln346_231_fu_12465_p3;
wire   [0:0] tmp_524_fu_12473_p3;
wire   [0:0] tmp_525_fu_12481_p3;
wire   [0:0] xor_ln895_190_fu_12489_p2;
wire   [0:0] and_ln895_135_fu_12495_p2;
wire   [0:0] xor_ln346_33_fu_12509_p2;
wire   [20:0] select_ln346_232_fu_12501_p3;
wire   [20:0] select_ln346_150_fu_12524_p3;
wire   [0:0] tmp_527_fu_12556_p3;
wire   [0:0] tmp_528_fu_12564_p3;
wire   [0:0] tmp_526_fu_12548_p3;
wire   [0:0] or_ln895_64_fu_12572_p2;
wire   [0:0] xor_ln895_191_fu_12578_p2;
wire   [0:0] and_ln896_65_fu_12590_p2;
wire   [0:0] xor_ln896_161_fu_12596_p2;
wire   [0:0] and_ln895_136_fu_12584_p2;
wire   [0:0] and_ln896_66_fu_12602_p2;
wire   [0:0] or_ln346_64_fu_12616_p2;
wire   [20:0] select_ln346_234_fu_12608_p3;
wire   [34:0] shl_ln1273_11_fu_12631_p3;
wire  signed [35:0] sext_ln1273_50_fu_12638_p1;
wire   [35:0] sub_ln1273_6_fu_12642_p2;
wire   [0:0] tmp_530_fu_12666_p3;
wire   [0:0] tmp_531_fu_12674_p3;
wire   [0:0] tmp_529_fu_12648_p3;
wire   [0:0] or_ln895_65_fu_12682_p2;
wire   [0:0] xor_ln895_192_fu_12688_p2;
wire   [0:0] and_ln896_67_fu_12700_p2;
wire   [0:0] xor_ln896_191_fu_12706_p2;
wire   [0:0] and_ln895_137_fu_12694_p2;
wire   [0:0] and_ln896_68_fu_12712_p2;
wire   [0:0] or_ln346_65_fu_12726_p2;
wire   [20:0] select_ln346_236_fu_12718_p3;
wire   [20:0] trunc_ln818_62_fu_12656_p4;
wire   [20:0] select_ln346_237_fu_12732_p3;
wire   [0:0] tmp_532_fu_12740_p3;
wire   [0:0] tmp_533_fu_12748_p3;
wire   [0:0] xor_ln895_193_fu_12756_p2;
wire   [0:0] and_ln895_138_fu_12762_p2;
wire   [0:0] xor_ln346_34_fu_12776_p2;
wire   [20:0] select_ln346_238_fu_12768_p3;
wire   [20:0] select_ln346_239_fu_12782_p3;
wire   [0:0] tmp_534_fu_12790_p3;
wire   [0:0] tmp_535_fu_12798_p3;
wire   [0:0] xor_ln895_194_fu_12806_p2;
wire   [0:0] and_ln895_139_fu_12812_p2;
wire   [0:0] xor_ln346_35_fu_12826_p2;
wire   [20:0] select_ln346_240_fu_12818_p3;
wire   [34:0] shl_ln1273_s_fu_12841_p3;
wire   [34:0] shl_ln1273_10_fu_12852_p3;
wire  signed [35:0] sext_ln810_fu_12848_p1;
wire   [35:0] sub_ln1273_7_fu_12863_p2;
wire   [0:0] tmp_537_fu_12887_p3;
wire   [0:0] tmp_538_fu_12895_p3;
wire   [0:0] tmp_536_fu_12869_p3;
wire   [0:0] or_ln895_66_fu_12903_p2;
wire   [0:0] xor_ln895_195_fu_12909_p2;
wire   [0:0] and_ln896_69_fu_12921_p2;
wire   [0:0] xor_ln896_192_fu_12927_p2;
wire   [0:0] and_ln895_140_fu_12915_p2;
wire   [0:0] and_ln896_70_fu_12933_p2;
wire   [0:0] or_ln346_66_fu_12947_p2;
wire   [20:0] select_ln346_242_fu_12939_p3;
wire   [20:0] trunc_ln818_63_fu_12877_p4;
wire   [20:0] select_ln346_243_fu_12953_p3;
wire   [0:0] tmp_539_fu_12961_p3;
wire   [0:0] tmp_540_fu_12969_p3;
wire   [0:0] xor_ln895_196_fu_12977_p2;
wire   [0:0] and_ln895_141_fu_12983_p2;
wire   [0:0] xor_ln346_36_fu_12997_p2;
wire   [20:0] select_ln346_244_fu_12989_p3;
wire  signed [35:0] sext_ln810_1_fu_12859_p1;
wire   [35:0] sub_ln1273_8_fu_13012_p2;
wire   [0:0] tmp_542_fu_13036_p3;
wire   [0:0] tmp_543_fu_13044_p3;
wire   [0:0] tmp_541_fu_13018_p3;
wire   [0:0] or_ln895_67_fu_13052_p2;
wire   [0:0] xor_ln895_197_fu_13058_p2;
wire   [0:0] and_ln896_71_fu_13070_p2;
wire   [0:0] xor_ln896_193_fu_13076_p2;
wire   [0:0] and_ln895_142_fu_13064_p2;
wire   [0:0] and_ln896_72_fu_13082_p2;
wire   [0:0] or_ln346_67_fu_13096_p2;
wire   [20:0] select_ln346_246_fu_13088_p3;
wire   [20:0] trunc_ln818_64_fu_13026_p4;
wire  signed [34:0] grp_fu_21654_p2;
wire   [0:0] tmp_349_fu_13134_p3;
wire   [20:0] zext_ln377_39_fu_13141_p1;
wire   [20:0] trunc_ln818_38_fu_13118_p4;
wire   [0:0] tmp_350_fu_13151_p3;
wire   [0:0] tmp_348_fu_13127_p3;
wire   [0:0] xor_ln896_96_fu_13159_p2;
wire   [0:0] xor_ln888_78_fu_13178_p2;
wire   [0:0] tmp_351_fu_13171_p3;
wire   [0:0] or_ln888_39_fu_13184_p2;
wire   [0:0] tmp_352_fu_13196_p3;
wire   [0:0] xor_ln890_39_fu_13203_p2;
wire   [0:0] or_ln890_39_fu_13209_p2;
wire   [0:0] and_ln378_39_fu_13165_p2;
wire   [0:0] xor_ln888_79_fu_13190_p2;
wire   [0:0] xor_ln895_126_fu_13227_p2;
wire   [0:0] tmp_347_fu_13111_p3;
wire   [0:0] or_ln895_39_fu_13233_p2;
wire   [0:0] xor_ln895_127_fu_13239_p2;
wire   [0:0] and_ln890_39_fu_13215_p2;
wire   [0:0] xor_ln896_97_fu_13251_p2;
wire   [0:0] and_ln891_39_fu_13221_p2;
wire   [0:0] or_ln896_39_fu_13257_p2;
wire   [0:0] xor_ln896_167_fu_13263_p2;
wire   [0:0] and_ln896_39_fu_13269_p2;
wire  signed [27:0] grp_fu_21666_p2;
wire   [13:0] trunc_ln818_39_fu_13288_p4;
wire   [0:0] tmp_359_fu_13308_p3;
wire   [14:0] zext_ln377_40_fu_13315_p1;
wire  signed [14:0] sext_ln365_2_fu_13297_p1;
wire   [0:0] tmp_360_fu_13325_p3;
wire   [0:0] tmp_358_fu_13301_p3;
wire   [0:0] xor_ln896_100_fu_13333_p2;
wire   [0:0] xor_ln888_80_fu_13352_p2;
wire   [0:0] tmp_361_fu_13345_p3;
wire   [0:0] or_ln888_40_fu_13358_p2;
wire   [0:0] tmp_362_fu_13370_p3;
wire   [0:0] xor_ln890_40_fu_13377_p2;
wire   [0:0] or_ln890_40_fu_13383_p2;
wire   [0:0] and_ln378_40_fu_13339_p2;
wire   [0:0] xor_ln888_81_fu_13364_p2;
wire   [0:0] xor_ln895_130_fu_13401_p2;
wire   [0:0] tmp_357_fu_13281_p3;
wire   [0:0] or_ln895_40_fu_13407_p2;
wire   [0:0] xor_ln895_131_fu_13413_p2;
wire   [0:0] and_ln890_40_fu_13389_p2;
wire   [0:0] xor_ln896_101_fu_13425_p2;
wire   [0:0] and_ln891_40_fu_13395_p2;
wire   [0:0] or_ln896_40_fu_13431_p2;
wire   [0:0] xor_ln896_168_fu_13437_p2;
wire   [0:0] and_ln896_40_fu_13443_p2;
wire  signed [34:0] grp_fu_21678_p2;
wire   [0:0] tmp_369_fu_13478_p3;
wire   [20:0] zext_ln377_41_fu_13485_p1;
wire   [20:0] trunc_ln818_40_fu_13462_p4;
wire   [20:0] add_ln377_41_fu_13489_p2;
wire   [0:0] tmp_370_fu_13495_p3;
wire   [0:0] tmp_368_fu_13471_p3;
wire   [0:0] xor_ln896_104_fu_13503_p2;
wire   [0:0] xor_ln888_82_fu_13522_p2;
wire   [0:0] tmp_371_fu_13515_p3;
wire   [0:0] or_ln888_41_fu_13528_p2;
wire   [0:0] tmp_372_fu_13540_p3;
wire   [0:0] xor_ln890_41_fu_13547_p2;
wire   [0:0] or_ln890_41_fu_13553_p2;
wire   [0:0] and_ln378_41_fu_13509_p2;
wire   [0:0] xor_ln888_83_fu_13534_p2;
wire   [0:0] xor_ln895_134_fu_13571_p2;
wire   [0:0] tmp_367_fu_13455_p3;
wire   [0:0] or_ln895_41_fu_13577_p2;
wire   [0:0] xor_ln895_135_fu_13583_p2;
wire   [0:0] and_ln890_41_fu_13559_p2;
wire   [0:0] xor_ln896_105_fu_13595_p2;
wire   [0:0] and_ln891_41_fu_13565_p2;
wire   [0:0] or_ln896_41_fu_13601_p2;
wire   [0:0] xor_ln896_169_fu_13607_p2;
wire   [0:0] and_ln895_101_fu_13589_p2;
wire   [0:0] and_ln896_41_fu_13613_p2;
wire   [0:0] or_ln346_41_fu_13619_p2;
wire   [20:0] select_ln346_164_fu_13625_p3;
wire  signed [28:0] grp_fu_21690_p2;
wire   [14:0] trunc_ln818_42_fu_13648_p4;
wire   [0:0] tmp_383_fu_13668_p3;
wire   [15:0] zext_ln377_43_fu_13675_p1;
wire  signed [15:0] sext_ln365_3_fu_13657_p1;
wire   [0:0] tmp_384_fu_13685_p3;
wire   [0:0] tmp_382_fu_13661_p3;
wire   [0:0] xor_ln896_109_fu_13693_p2;
wire   [0:0] xor_ln888_86_fu_13712_p2;
wire   [0:0] tmp_385_fu_13705_p3;
wire   [0:0] or_ln888_43_fu_13718_p2;
wire   [0:0] tmp_386_fu_13730_p3;
wire   [0:0] xor_ln890_43_fu_13737_p2;
wire   [0:0] or_ln890_43_fu_13743_p2;
wire   [0:0] and_ln378_43_fu_13699_p2;
wire   [0:0] xor_ln888_87_fu_13724_p2;
wire   [0:0] xor_ln895_139_fu_13761_p2;
wire   [0:0] tmp_381_fu_13641_p3;
wire   [0:0] or_ln895_43_fu_13767_p2;
wire   [0:0] xor_ln895_140_fu_13773_p2;
wire   [0:0] and_ln890_43_fu_13749_p2;
wire   [0:0] xor_ln896_110_fu_13785_p2;
wire   [0:0] and_ln891_43_fu_13755_p2;
wire   [0:0] or_ln896_43_fu_13791_p2;
wire   [0:0] xor_ln896_171_fu_13797_p2;
wire   [0:0] and_ln896_43_fu_13803_p2;
wire  signed [33:0] grp_fu_21702_p2;
wire   [19:0] trunc_ln818_44_fu_13822_p4;
wire   [0:0] tmp_397_fu_13842_p3;
wire   [20:0] zext_ln377_45_fu_13849_p1;
wire  signed [20:0] sext_ln818_1_fu_13831_p1;
wire   [20:0] add_ln377_45_fu_13853_p2;
wire   [0:0] tmp_398_fu_13859_p3;
wire   [0:0] tmp_396_fu_13835_p3;
wire   [0:0] xor_ln896_114_fu_13867_p2;
wire   [0:0] xor_ln888_90_fu_13886_p2;
wire   [0:0] tmp_399_fu_13879_p3;
wire   [0:0] or_ln888_45_fu_13892_p2;
wire   [0:0] tmp_400_fu_13904_p3;
wire   [0:0] xor_ln890_45_fu_13911_p2;
wire   [0:0] or_ln890_45_fu_13917_p2;
wire   [0:0] and_ln378_45_fu_13873_p2;
wire   [0:0] xor_ln888_91_fu_13898_p2;
wire   [0:0] xor_ln895_144_fu_13935_p2;
wire   [0:0] tmp_395_fu_13815_p3;
wire   [0:0] or_ln895_45_fu_13941_p2;
wire   [0:0] xor_ln895_145_fu_13947_p2;
wire   [0:0] and_ln890_45_fu_13923_p2;
wire   [0:0] xor_ln896_115_fu_13959_p2;
wire   [0:0] and_ln891_45_fu_13929_p2;
wire   [0:0] or_ln896_45_fu_13965_p2;
wire   [0:0] xor_ln896_173_fu_13971_p2;
wire   [0:0] and_ln895_107_fu_13953_p2;
wire   [0:0] and_ln896_45_fu_13977_p2;
wire   [0:0] or_ln346_45_fu_13983_p2;
wire   [20:0] select_ln346_176_fu_13989_p3;
wire  signed [29:0] grp_fu_21721_p2;
wire   [15:0] trunc_ln818_47_fu_14019_p4;
wire   [0:0] tmp_415_fu_14039_p3;
wire   [16:0] zext_ln377_48_fu_14046_p1;
wire  signed [16:0] sext_ln365_4_fu_14028_p1;
wire   [0:0] tmp_416_fu_14056_p3;
wire   [0:0] tmp_414_fu_14032_p3;
wire   [0:0] xor_ln896_120_fu_14064_p2;
wire   [0:0] xor_ln888_96_fu_14083_p2;
wire   [0:0] tmp_417_fu_14076_p3;
wire   [0:0] or_ln888_48_fu_14089_p2;
wire   [0:0] tmp_418_fu_14101_p3;
wire   [0:0] xor_ln890_48_fu_14108_p2;
wire   [0:0] or_ln890_48_fu_14114_p2;
wire   [0:0] and_ln378_48_fu_14070_p2;
wire   [0:0] xor_ln888_97_fu_14095_p2;
wire   [0:0] xor_ln895_150_fu_14132_p2;
wire   [0:0] tmp_413_fu_14012_p3;
wire   [0:0] or_ln895_48_fu_14138_p2;
wire   [0:0] xor_ln895_151_fu_14144_p2;
wire   [0:0] and_ln890_48_fu_14120_p2;
wire   [0:0] xor_ln896_121_fu_14156_p2;
wire   [0:0] and_ln891_48_fu_14126_p2;
wire   [0:0] or_ln896_48_fu_14162_p2;
wire   [0:0] xor_ln896_176_fu_14168_p2;
wire   [0:0] and_ln896_48_fu_14174_p2;
wire  signed [34:0] grp_fu_21740_p2;
wire   [0:0] tmp_453_fu_14216_p3;
wire   [20:0] zext_ln377_53_fu_14223_p1;
wire   [20:0] trunc_ln818_52_fu_14200_p4;
wire   [20:0] add_ln377_53_fu_14227_p2;
wire   [0:0] tmp_454_fu_14233_p3;
wire   [0:0] tmp_452_fu_14209_p3;
wire   [0:0] xor_ln896_134_fu_14241_p2;
wire   [0:0] xor_ln888_106_fu_14260_p2;
wire   [0:0] tmp_455_fu_14253_p3;
wire   [0:0] or_ln888_53_fu_14266_p2;
wire   [0:0] tmp_456_fu_14278_p3;
wire   [0:0] xor_ln890_53_fu_14285_p2;
wire   [0:0] or_ln890_53_fu_14291_p2;
wire   [0:0] and_ln378_53_fu_14247_p2;
wire   [0:0] xor_ln888_107_fu_14272_p2;
wire   [0:0] xor_ln895_164_fu_14309_p2;
wire   [0:0] tmp_451_fu_14193_p3;
wire   [0:0] or_ln895_53_fu_14315_p2;
wire   [0:0] xor_ln895_165_fu_14321_p2;
wire   [0:0] and_ln890_53_fu_14297_p2;
wire   [0:0] xor_ln896_135_fu_14333_p2;
wire   [0:0] and_ln891_53_fu_14303_p2;
wire   [0:0] or_ln896_53_fu_14339_p2;
wire   [0:0] xor_ln896_181_fu_14345_p2;
wire   [0:0] and_ln895_119_fu_14327_p2;
wire   [0:0] and_ln896_53_fu_14351_p2;
wire   [0:0] or_ln346_53_fu_14357_p2;
wire   [20:0] select_ln346_200_fu_14363_p3;
wire  signed [28:0] grp_fu_21752_p2;
wire   [14:0] trunc_ln818_54_fu_14386_p4;
wire   [0:0] tmp_467_fu_14406_p3;
wire   [15:0] zext_ln377_55_fu_14413_p1;
wire  signed [15:0] sext_ln365_6_fu_14395_p1;
wire   [0:0] tmp_468_fu_14423_p3;
wire   [0:0] tmp_466_fu_14399_p3;
wire   [0:0] xor_ln896_139_fu_14431_p2;
wire   [0:0] xor_ln888_110_fu_14450_p2;
wire   [0:0] tmp_469_fu_14443_p3;
wire   [0:0] or_ln888_55_fu_14456_p2;
wire   [0:0] tmp_470_fu_14468_p3;
wire   [0:0] xor_ln890_55_fu_14475_p2;
wire   [0:0] or_ln890_55_fu_14481_p2;
wire   [0:0] and_ln378_55_fu_14437_p2;
wire   [0:0] xor_ln888_111_fu_14462_p2;
wire   [0:0] xor_ln895_169_fu_14499_p2;
wire   [0:0] tmp_465_fu_14379_p3;
wire   [0:0] or_ln895_55_fu_14505_p2;
wire   [0:0] xor_ln895_170_fu_14511_p2;
wire   [0:0] and_ln890_55_fu_14487_p2;
wire   [0:0] xor_ln896_140_fu_14523_p2;
wire   [0:0] and_ln891_55_fu_14493_p2;
wire   [0:0] or_ln896_55_fu_14529_p2;
wire   [0:0] xor_ln896_183_fu_14535_p2;
wire   [0:0] and_ln896_55_fu_14541_p2;
wire  signed [33:0] grp_fu_21764_p2;
wire   [19:0] trunc_ln818_56_fu_14560_p4;
wire   [0:0] tmp_481_fu_14580_p3;
wire   [20:0] zext_ln377_57_fu_14587_p1;
wire  signed [20:0] sext_ln818_2_fu_14569_p1;
wire   [20:0] add_ln377_57_fu_14591_p2;
wire   [0:0] tmp_482_fu_14597_p3;
wire   [0:0] tmp_480_fu_14573_p3;
wire   [0:0] xor_ln896_144_fu_14605_p2;
wire   [0:0] xor_ln888_114_fu_14624_p2;
wire   [0:0] tmp_483_fu_14617_p3;
wire   [0:0] or_ln888_57_fu_14630_p2;
wire   [0:0] tmp_484_fu_14642_p3;
wire   [0:0] xor_ln890_57_fu_14649_p2;
wire   [0:0] or_ln890_57_fu_14655_p2;
wire   [0:0] and_ln378_57_fu_14611_p2;
wire   [0:0] xor_ln888_115_fu_14636_p2;
wire   [0:0] xor_ln895_174_fu_14673_p2;
wire   [0:0] tmp_479_fu_14553_p3;
wire   [0:0] or_ln895_57_fu_14679_p2;
wire   [0:0] xor_ln895_175_fu_14685_p2;
wire   [0:0] and_ln890_57_fu_14661_p2;
wire   [0:0] xor_ln896_145_fu_14697_p2;
wire   [0:0] and_ln891_57_fu_14667_p2;
wire   [0:0] or_ln896_57_fu_14703_p2;
wire   [0:0] xor_ln896_185_fu_14709_p2;
wire   [0:0] and_ln895_125_fu_14691_p2;
wire   [0:0] and_ln896_57_fu_14715_p2;
wire   [0:0] or_ln346_57_fu_14721_p2;
wire   [20:0] select_ln346_212_fu_14727_p3;
wire  signed [29:0] grp_fu_21783_p2;
wire   [15:0] trunc_ln818_59_fu_14757_p4;
wire   [0:0] tmp_499_fu_14777_p3;
wire   [16:0] zext_ln377_60_fu_14784_p1;
wire  signed [16:0] sext_ln365_7_fu_14766_p1;
wire   [0:0] tmp_500_fu_14794_p3;
wire   [0:0] tmp_498_fu_14770_p3;
wire   [0:0] xor_ln896_150_fu_14802_p2;
wire   [0:0] xor_ln888_120_fu_14821_p2;
wire   [0:0] tmp_501_fu_14814_p3;
wire   [0:0] or_ln888_60_fu_14827_p2;
wire   [0:0] tmp_502_fu_14839_p3;
wire   [0:0] xor_ln890_60_fu_14846_p2;
wire   [0:0] or_ln890_60_fu_14852_p2;
wire   [0:0] and_ln378_60_fu_14808_p2;
wire   [0:0] xor_ln888_121_fu_14833_p2;
wire   [0:0] xor_ln895_180_fu_14870_p2;
wire   [0:0] tmp_497_fu_14750_p3;
wire   [0:0] or_ln895_60_fu_14876_p2;
wire   [0:0] xor_ln895_181_fu_14882_p2;
wire   [0:0] and_ln890_60_fu_14858_p2;
wire   [0:0] xor_ln896_151_fu_14894_p2;
wire   [0:0] and_ln891_60_fu_14864_p2;
wire   [0:0] or_ln896_60_fu_14900_p2;
wire   [0:0] xor_ln896_188_fu_14906_p2;
wire   [0:0] and_ln896_60_fu_14912_p2;
wire   [20:0] select_ln346_152_fu_14931_p3;
wire   [20:0] select_ln346_153_fu_14938_p3;
wire   [0:0] tmp_353_fu_14944_p3;
wire   [0:0] tmp_354_fu_14952_p3;
wire   [0:0] xor_ln895_128_fu_14960_p2;
wire   [0:0] and_ln895_96_fu_14966_p2;
wire   [0:0] xor_ln346_18_fu_14980_p2;
wire   [20:0] select_ln346_154_fu_14972_p3;
wire   [20:0] select_ln346_155_fu_14986_p3;
wire   [0:0] tmp_355_fu_14994_p3;
wire   [0:0] tmp_356_fu_15002_p3;
wire   [0:0] xor_ln895_129_fu_15010_p2;
wire   [0:0] and_ln895_97_fu_15016_p2;
wire   [0:0] xor_ln346_19_fu_15030_p2;
wire   [20:0] select_ln346_156_fu_15022_p3;
wire   [20:0] select_ln346_158_fu_15048_p3;
wire  signed [20:0] sext_ln856_2_fu_15045_p1;
wire   [20:0] select_ln346_159_fu_15055_p3;
wire   [0:0] tmp_363_fu_15062_p3;
wire   [0:0] tmp_364_fu_15070_p3;
wire   [0:0] xor_ln895_132_fu_15078_p2;
wire   [0:0] and_ln895_99_fu_15084_p2;
wire   [0:0] xor_ln346_20_fu_15098_p2;
wire   [20:0] select_ln346_160_fu_15090_p3;
wire   [20:0] select_ln346_161_fu_15104_p3;
wire   [0:0] tmp_365_fu_15112_p3;
wire   [0:0] tmp_366_fu_15120_p3;
wire   [0:0] xor_ln895_133_fu_15128_p2;
wire   [0:0] and_ln895_100_fu_15134_p2;
wire   [0:0] xor_ln346_21_fu_15148_p2;
wire   [20:0] select_ln346_162_fu_15140_p3;
wire  signed [34:0] shl_ln838_32_fu_15163_p3;
wire  signed [34:0] grp_fu_21802_p2;
wire  signed [35:0] sext_ln813_110_fu_15170_p1;
wire  signed [35:0] sext_ln1347_46_fu_15174_p1;
wire   [35:0] add_ln1347_51_fu_15177_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_27_fu_15183_p2;
wire   [0:0] tmp_375_fu_15214_p3;
wire   [20:0] zext_ln377_42_fu_15221_p1;
wire   [20:0] trunc_ln818_41_fu_15196_p4;
wire   [0:0] tmp_376_fu_15231_p3;
wire   [0:0] xor_ln888_84_fu_15253_p2;
wire   [0:0] or_ln888_42_fu_15259_p2;
wire   [0:0] tmp_378_fu_15271_p3;
wire   [0:0] xor_ln890_42_fu_15279_p2;
wire   [0:0] or_ln890_42_fu_15285_p2;
wire   [0:0] xor_ln888_85_fu_15265_p2;
wire   [0:0] xor_ln895_136_fu_15297_p2;
wire   [0:0] or_ln895_42_fu_15303_p2;
wire   [0:0] xor_ln895_137_fu_15309_p2;
wire   [0:0] and_ln890_42_fu_15291_p2;
wire   [0:0] xor_ln896_107_fu_15321_p2;
wire   [20:0] select_ln346_170_fu_15336_p3;
wire  signed [20:0] sext_ln856_3_fu_15333_p1;
wire   [20:0] select_ln346_171_fu_15343_p3;
wire  signed [34:0] shl_ln838_33_fu_15350_p3;
wire  signed [27:0] grp_fu_21810_p2;
wire  signed [35:0] sext_ln813_111_fu_15358_p1;
wire  signed [35:0] sext_ln1347_47_fu_15362_p1;
wire  signed [34:0] sext_ln1347_48_fu_15365_p1;
wire   [35:0] add_ln1347_52_fu_15368_p2;
wire   [34:0] add_ln810_28_fu_15374_p2;
wire   [0:0] tmp_389_fu_15406_p3;
wire   [20:0] zext_ln377_44_fu_15413_p1;
wire   [20:0] trunc_ln818_43_fu_15388_p4;
wire   [0:0] tmp_390_fu_15423_p3;
wire   [0:0] xor_ln888_88_fu_15445_p2;
wire   [0:0] or_ln888_44_fu_15451_p2;
wire   [0:0] tmp_392_fu_15463_p3;
wire   [0:0] xor_ln890_44_fu_15471_p2;
wire   [0:0] or_ln890_44_fu_15477_p2;
wire   [0:0] xor_ln888_89_fu_15457_p2;
wire   [0:0] xor_ln895_141_fu_15489_p2;
wire   [0:0] or_ln895_44_fu_15495_p2;
wire   [0:0] xor_ln895_142_fu_15501_p2;
wire   [0:0] and_ln890_44_fu_15483_p2;
wire   [0:0] xor_ln896_112_fu_15513_p2;
wire  signed [34:0] shl_ln838_34_fu_15525_p3;
wire  signed [35:0] sext_ln813_112_fu_15532_p1;
wire  signed [35:0] sext_ln1347_49_fu_15536_p1;
wire   [35:0] add_ln1347_53_fu_15539_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_29_fu_15545_p2;
wire   [20:0] zext_ln377_46_fu_15576_p1;
wire   [20:0] trunc_ln818_45_fu_15558_p4;
wire   [20:0] add_ln377_46_fu_15579_p2;
wire   [0:0] tmp_404_fu_15585_p3;
wire   [0:0] tmp_402_fu_15568_p3;
wire   [0:0] xor_ln896_116_fu_15593_p2;
wire   [0:0] xor_ln888_92_fu_15613_p2;
wire   [0:0] tmp_405_fu_15605_p3;
wire   [0:0] or_ln888_46_fu_15619_p2;
wire   [0:0] tmp_406_fu_15631_p3;
wire   [0:0] xor_ln890_46_fu_15639_p2;
wire   [0:0] or_ln890_46_fu_15645_p2;
wire   [0:0] and_ln378_46_fu_15599_p2;
wire   [0:0] xor_ln888_93_fu_15625_p2;
wire   [0:0] xor_ln895_146_fu_15663_p2;
wire   [0:0] tmp_401_fu_15550_p3;
wire   [0:0] or_ln895_46_fu_15669_p2;
wire   [0:0] xor_ln895_147_fu_15675_p2;
wire   [0:0] and_ln890_46_fu_15651_p2;
wire   [0:0] xor_ln896_117_fu_15687_p2;
wire   [0:0] and_ln891_46_fu_15657_p2;
wire   [0:0] or_ln896_46_fu_15693_p2;
wire   [0:0] xor_ln896_174_fu_15699_p2;
wire   [0:0] and_ln895_108_fu_15681_p2;
wire   [0:0] and_ln896_46_fu_15705_p2;
wire   [0:0] or_ln346_46_fu_15711_p2;
wire   [20:0] select_ln346_178_fu_15717_p3;
wire   [20:0] select_ln346_182_fu_15743_p3;
wire  signed [20:0] sext_ln856_4_fu_15740_p1;
wire   [20:0] select_ln346_183_fu_15750_p3;
wire  signed [34:0] shl_ln838_36_fu_15757_p3;
wire  signed [35:0] sext_ln813_114_fu_15765_p1;
wire  signed [35:0] sext_ln1347_51_fu_15769_p1;
wire  signed [34:0] sext_ln1347_52_fu_15772_p1;
wire   [35:0] add_ln1347_55_fu_15775_p2;
wire   [34:0] add_ln810_31_fu_15781_p2;
wire   [20:0] zext_ln377_49_fu_15813_p1;
wire   [20:0] trunc_ln818_48_fu_15795_p4;
wire   [20:0] add_ln377_49_fu_15816_p2;
wire   [0:0] tmp_422_fu_15822_p3;
wire   [0:0] tmp_420_fu_15805_p3;
wire   [0:0] xor_ln896_122_fu_15830_p2;
wire   [0:0] xor_ln888_98_fu_15850_p2;
wire   [0:0] tmp_423_fu_15842_p3;
wire   [0:0] or_ln888_49_fu_15856_p2;
wire   [0:0] tmp_424_fu_15868_p3;
wire   [0:0] xor_ln890_49_fu_15876_p2;
wire   [0:0] or_ln890_49_fu_15882_p2;
wire   [0:0] and_ln378_49_fu_15836_p2;
wire   [0:0] xor_ln888_99_fu_15862_p2;
wire   [0:0] xor_ln895_152_fu_15900_p2;
wire   [0:0] tmp_419_fu_15787_p3;
wire   [0:0] or_ln895_49_fu_15906_p2;
wire   [0:0] xor_ln895_153_fu_15912_p2;
wire   [0:0] and_ln890_49_fu_15888_p2;
wire   [0:0] xor_ln896_123_fu_15924_p2;
wire   [0:0] and_ln891_49_fu_15894_p2;
wire   [0:0] or_ln896_49_fu_15930_p2;
wire   [0:0] xor_ln896_177_fu_15936_p2;
wire   [0:0] and_ln895_111_fu_15918_p2;
wire   [0:0] and_ln896_49_fu_15942_p2;
wire   [0:0] or_ln346_49_fu_15948_p2;
wire   [20:0] select_ln346_184_fu_15954_p3;
wire  signed [34:0] grp_fu_21833_p2;
wire   [0:0] tmp_433_fu_16000_p3;
wire   [20:0] zext_ln377_51_fu_16007_p1;
wire   [20:0] trunc_ln818_50_fu_15984_p4;
wire   [0:0] tmp_434_fu_16017_p3;
wire   [0:0] tmp_432_fu_15993_p3;
wire   [0:0] xor_ln896_126_fu_16025_p2;
wire   [0:0] xor_ln888_102_fu_16044_p2;
wire   [0:0] tmp_435_fu_16037_p3;
wire   [0:0] or_ln888_51_fu_16050_p2;
wire   [0:0] tmp_436_fu_16062_p3;
wire   [0:0] xor_ln890_51_fu_16069_p2;
wire   [0:0] or_ln890_51_fu_16075_p2;
wire   [0:0] and_ln378_51_fu_16031_p2;
wire   [0:0] xor_ln888_103_fu_16056_p2;
wire   [0:0] xor_ln895_156_fu_16093_p2;
wire   [0:0] tmp_431_fu_15977_p3;
wire   [0:0] or_ln895_51_fu_16099_p2;
wire   [0:0] xor_ln895_157_fu_16105_p2;
wire   [0:0] and_ln890_51_fu_16081_p2;
wire   [0:0] xor_ln896_127_fu_16117_p2;
wire   [0:0] and_ln891_51_fu_16087_p2;
wire   [0:0] or_ln896_51_fu_16123_p2;
wire   [0:0] xor_ln896_179_fu_16129_p2;
wire   [0:0] and_ln896_51_fu_16135_p2;
wire  signed [27:0] grp_fu_21844_p2;
wire   [13:0] trunc_ln818_51_fu_16154_p4;
wire   [0:0] tmp_443_fu_16174_p3;
wire   [14:0] zext_ln377_52_fu_16181_p1;
wire  signed [14:0] sext_ln365_5_fu_16163_p1;
wire   [0:0] tmp_444_fu_16191_p3;
wire   [0:0] tmp_442_fu_16167_p3;
wire   [0:0] xor_ln896_130_fu_16199_p2;
wire   [0:0] xor_ln888_104_fu_16218_p2;
wire   [0:0] tmp_445_fu_16211_p3;
wire   [0:0] or_ln888_52_fu_16224_p2;
wire   [0:0] tmp_446_fu_16236_p3;
wire   [0:0] xor_ln890_52_fu_16243_p2;
wire   [0:0] or_ln890_52_fu_16249_p2;
wire   [0:0] and_ln378_52_fu_16205_p2;
wire   [0:0] xor_ln888_105_fu_16230_p2;
wire   [0:0] xor_ln895_160_fu_16267_p2;
wire   [0:0] tmp_441_fu_16147_p3;
wire   [0:0] or_ln895_52_fu_16273_p2;
wire   [0:0] xor_ln895_161_fu_16279_p2;
wire   [0:0] and_ln890_52_fu_16255_p2;
wire   [0:0] xor_ln896_131_fu_16291_p2;
wire   [0:0] and_ln891_52_fu_16261_p2;
wire   [0:0] or_ln896_52_fu_16297_p2;
wire   [0:0] xor_ln896_180_fu_16303_p2;
wire   [0:0] and_ln896_52_fu_16309_p2;
wire  signed [34:0] shl_ln838_38_fu_16321_p3;
wire  signed [34:0] grp_fu_21855_p2;
wire  signed [35:0] sext_ln813_116_fu_16328_p1;
wire  signed [35:0] sext_ln1347_55_fu_16332_p1;
wire   [35:0] add_ln1347_57_fu_16335_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_33_fu_16341_p2;
wire   [0:0] tmp_459_fu_16372_p3;
wire   [20:0] zext_ln377_54_fu_16379_p1;
wire   [20:0] trunc_ln818_53_fu_16354_p4;
wire   [0:0] tmp_460_fu_16389_p3;
wire   [0:0] xor_ln888_108_fu_16411_p2;
wire   [0:0] or_ln888_54_fu_16417_p2;
wire   [0:0] tmp_462_fu_16429_p3;
wire   [0:0] xor_ln890_54_fu_16437_p2;
wire   [0:0] or_ln890_54_fu_16443_p2;
wire   [0:0] xor_ln888_109_fu_16423_p2;
wire   [0:0] xor_ln895_166_fu_16455_p2;
wire   [0:0] or_ln895_54_fu_16461_p2;
wire   [0:0] xor_ln895_167_fu_16467_p2;
wire   [0:0] and_ln890_54_fu_16449_p2;
wire   [0:0] xor_ln896_137_fu_16479_p2;
wire   [20:0] select_ln346_206_fu_16494_p3;
wire  signed [20:0] sext_ln856_6_fu_16491_p1;
wire   [20:0] select_ln346_207_fu_16501_p3;
wire  signed [34:0] shl_ln838_39_fu_16508_p3;
wire  signed [27:0] grp_fu_21863_p2;
wire  signed [35:0] sext_ln813_117_fu_16516_p1;
wire  signed [35:0] sext_ln1347_56_fu_16520_p1;
wire  signed [34:0] sext_ln1347_57_fu_16523_p1;
wire   [35:0] add_ln1347_58_fu_16526_p2;
wire   [34:0] add_ln810_34_fu_16532_p2;
wire   [0:0] tmp_473_fu_16564_p3;
wire   [20:0] zext_ln377_56_fu_16571_p1;
wire   [20:0] trunc_ln818_55_fu_16546_p4;
wire   [0:0] tmp_474_fu_16581_p3;
wire   [0:0] xor_ln888_112_fu_16603_p2;
wire   [0:0] or_ln888_56_fu_16609_p2;
wire   [0:0] tmp_476_fu_16621_p3;
wire   [0:0] xor_ln890_56_fu_16629_p2;
wire   [0:0] or_ln890_56_fu_16635_p2;
wire   [0:0] xor_ln888_113_fu_16615_p2;
wire   [0:0] xor_ln895_171_fu_16647_p2;
wire   [0:0] or_ln895_56_fu_16653_p2;
wire   [0:0] xor_ln895_172_fu_16659_p2;
wire   [0:0] and_ln890_56_fu_16641_p2;
wire   [0:0] xor_ln896_142_fu_16671_p2;
wire  signed [34:0] shl_ln838_40_fu_16683_p3;
wire  signed [35:0] sext_ln813_118_fu_16690_p1;
wire  signed [35:0] sext_ln1347_58_fu_16694_p1;
wire   [35:0] add_ln1347_59_fu_16697_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_35_fu_16703_p2;
wire   [20:0] zext_ln377_58_fu_16734_p1;
wire   [20:0] trunc_ln818_57_fu_16716_p4;
wire   [20:0] add_ln377_58_fu_16737_p2;
wire   [0:0] tmp_488_fu_16743_p3;
wire   [0:0] tmp_486_fu_16726_p3;
wire   [0:0] xor_ln896_146_fu_16751_p2;
wire   [0:0] xor_ln888_116_fu_16771_p2;
wire   [0:0] tmp_489_fu_16763_p3;
wire   [0:0] or_ln888_58_fu_16777_p2;
wire   [0:0] tmp_490_fu_16789_p3;
wire   [0:0] xor_ln890_58_fu_16797_p2;
wire   [0:0] or_ln890_58_fu_16803_p2;
wire   [0:0] and_ln378_58_fu_16757_p2;
wire   [0:0] xor_ln888_117_fu_16783_p2;
wire   [0:0] xor_ln895_176_fu_16821_p2;
wire   [0:0] tmp_485_fu_16708_p3;
wire   [0:0] or_ln895_58_fu_16827_p2;
wire   [0:0] xor_ln895_177_fu_16833_p2;
wire   [0:0] and_ln890_58_fu_16809_p2;
wire   [0:0] xor_ln896_147_fu_16845_p2;
wire   [0:0] and_ln891_58_fu_16815_p2;
wire   [0:0] or_ln896_58_fu_16851_p2;
wire   [0:0] xor_ln896_186_fu_16857_p2;
wire   [0:0] and_ln895_126_fu_16839_p2;
wire   [0:0] and_ln896_58_fu_16863_p2;
wire   [0:0] or_ln346_58_fu_16869_p2;
wire   [20:0] select_ln346_214_fu_16875_p3;
wire   [20:0] select_ln346_218_fu_16901_p3;
wire  signed [20:0] sext_ln856_7_fu_16898_p1;
wire   [20:0] select_ln346_219_fu_16908_p3;
wire  signed [34:0] shl_ln838_42_fu_16915_p3;
wire  signed [35:0] sext_ln813_120_fu_16923_p1;
wire  signed [35:0] sext_ln1347_60_fu_16927_p1;
wire  signed [34:0] sext_ln1347_61_fu_16930_p1;
wire   [35:0] add_ln1347_61_fu_16933_p2;
wire   [34:0] add_ln810_37_fu_16939_p2;
wire   [20:0] zext_ln377_61_fu_16971_p1;
wire   [20:0] trunc_ln818_60_fu_16953_p4;
wire   [20:0] add_ln377_61_fu_16974_p2;
wire   [0:0] tmp_506_fu_16980_p3;
wire   [0:0] tmp_504_fu_16963_p3;
wire   [0:0] xor_ln896_152_fu_16988_p2;
wire   [0:0] xor_ln888_122_fu_17008_p2;
wire   [0:0] tmp_507_fu_17000_p3;
wire   [0:0] or_ln888_61_fu_17014_p2;
wire   [0:0] tmp_508_fu_17026_p3;
wire   [0:0] xor_ln890_61_fu_17034_p2;
wire   [0:0] or_ln890_61_fu_17040_p2;
wire   [0:0] and_ln378_61_fu_16994_p2;
wire   [0:0] xor_ln888_123_fu_17020_p2;
wire   [0:0] xor_ln895_182_fu_17058_p2;
wire   [0:0] tmp_503_fu_16945_p3;
wire   [0:0] or_ln895_61_fu_17064_p2;
wire   [0:0] xor_ln895_183_fu_17070_p2;
wire   [0:0] and_ln890_61_fu_17046_p2;
wire   [0:0] xor_ln896_153_fu_17082_p2;
wire   [0:0] and_ln891_61_fu_17052_p2;
wire   [0:0] or_ln896_61_fu_17088_p2;
wire   [0:0] xor_ln896_189_fu_17094_p2;
wire   [0:0] and_ln895_129_fu_17076_p2;
wire   [0:0] and_ln896_61_fu_17100_p2;
wire   [0:0] or_ln346_61_fu_17106_p2;
wire   [20:0] select_ln346_220_fu_17112_p3;
wire   [0:0] and_ln378_42_fu_17135_p2;
wire   [0:0] and_ln891_42_fu_17139_p2;
wire   [0:0] xor_ln896_170_fu_17144_p2;
wire   [0:0] and_ln896_42_fu_17149_p2;
wire   [0:0] or_ln346_42_fu_17161_p2;
wire   [20:0] select_ln346_166_fu_17154_p3;
wire   [20:0] select_ln346_167_fu_17166_p3;
wire   [0:0] tmp_379_fu_17173_p3;
wire   [0:0] tmp_380_fu_17181_p3;
wire   [0:0] xor_ln895_138_fu_17189_p2;
wire   [0:0] and_ln895_103_fu_17195_p2;
wire   [0:0] xor_ln346_22_fu_17209_p2;
wire   [20:0] select_ln346_168_fu_17201_p3;
wire   [0:0] and_ln378_44_fu_17223_p2;
wire   [0:0] and_ln891_44_fu_17227_p2;
wire   [0:0] xor_ln896_172_fu_17232_p2;
wire   [0:0] and_ln896_44_fu_17237_p2;
wire   [0:0] or_ln346_44_fu_17249_p2;
wire   [20:0] select_ln346_172_fu_17242_p3;
wire   [20:0] select_ln346_173_fu_17254_p3;
wire   [0:0] tmp_393_fu_17261_p3;
wire   [0:0] tmp_394_fu_17269_p3;
wire   [0:0] xor_ln895_143_fu_17277_p2;
wire   [0:0] and_ln895_106_fu_17283_p2;
wire   [0:0] xor_ln346_23_fu_17297_p2;
wire   [20:0] select_ln346_174_fu_17289_p3;
wire  signed [34:0] shl_ln838_35_fu_17311_p3;
wire  signed [35:0] sext_ln813_113_fu_17318_p1;
wire  signed [35:0] sext_ln1347_50_fu_17322_p1;
wire   [35:0] add_ln1347_54_fu_17325_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_30_fu_17331_p2;
wire   [20:0] zext_ln377_47_fu_17362_p1;
wire   [20:0] trunc_ln818_46_fu_17344_p4;
wire   [20:0] add_ln377_47_fu_17365_p2;
wire   [0:0] tmp_410_fu_17371_p3;
wire   [0:0] tmp_408_fu_17354_p3;
wire   [0:0] xor_ln896_118_fu_17379_p2;
wire   [0:0] xor_ln888_94_fu_17399_p2;
wire   [0:0] tmp_411_fu_17391_p3;
wire   [0:0] or_ln888_47_fu_17405_p2;
wire   [0:0] tmp_412_fu_17417_p3;
wire   [0:0] xor_ln890_47_fu_17425_p2;
wire   [0:0] or_ln890_47_fu_17431_p2;
wire   [0:0] and_ln378_47_fu_17385_p2;
wire   [0:0] xor_ln888_95_fu_17411_p2;
wire   [0:0] xor_ln895_148_fu_17449_p2;
wire   [0:0] tmp_407_fu_17336_p3;
wire   [0:0] or_ln895_47_fu_17455_p2;
wire   [0:0] xor_ln895_149_fu_17461_p2;
wire   [0:0] and_ln890_47_fu_17437_p2;
wire   [0:0] xor_ln896_119_fu_17473_p2;
wire   [0:0] and_ln891_47_fu_17443_p2;
wire   [0:0] or_ln896_47_fu_17479_p2;
wire   [0:0] xor_ln896_175_fu_17485_p2;
wire   [0:0] and_ln895_109_fu_17467_p2;
wire   [0:0] and_ln896_47_fu_17491_p2;
wire   [0:0] or_ln346_47_fu_17505_p2;
wire   [20:0] select_ln346_180_fu_17497_p3;
wire  signed [34:0] shl_ln838_37_fu_17519_p3;
wire  signed [35:0] sext_ln813_115_fu_17526_p1;
wire  signed [35:0] sext_ln1347_53_fu_17530_p1;
wire  signed [34:0] sext_ln1347_54_fu_17533_p1;
wire   [35:0] add_ln1347_56_fu_17536_p2;
wire   [34:0] add_ln810_32_fu_17542_p2;
wire   [20:0] zext_ln377_50_fu_17574_p1;
wire   [20:0] trunc_ln818_49_fu_17556_p4;
wire   [20:0] add_ln377_50_fu_17577_p2;
wire   [0:0] tmp_428_fu_17583_p3;
wire   [0:0] tmp_426_fu_17566_p3;
wire   [0:0] xor_ln896_124_fu_17591_p2;
wire   [0:0] xor_ln888_100_fu_17611_p2;
wire   [0:0] tmp_429_fu_17603_p3;
wire   [0:0] or_ln888_50_fu_17617_p2;
wire   [0:0] tmp_430_fu_17629_p3;
wire   [0:0] xor_ln890_50_fu_17637_p2;
wire   [0:0] or_ln890_50_fu_17643_p2;
wire   [0:0] and_ln378_50_fu_17597_p2;
wire   [0:0] xor_ln888_101_fu_17623_p2;
wire   [0:0] xor_ln895_154_fu_17661_p2;
wire   [0:0] tmp_425_fu_17548_p3;
wire   [0:0] or_ln895_50_fu_17667_p2;
wire   [0:0] xor_ln895_155_fu_17673_p2;
wire   [0:0] and_ln890_50_fu_17649_p2;
wire   [0:0] xor_ln896_125_fu_17685_p2;
wire   [0:0] and_ln891_50_fu_17655_p2;
wire   [0:0] or_ln896_50_fu_17691_p2;
wire   [0:0] xor_ln896_178_fu_17697_p2;
wire   [0:0] and_ln895_112_fu_17679_p2;
wire   [0:0] and_ln896_50_fu_17703_p2;
wire   [0:0] or_ln346_50_fu_17717_p2;
wire   [20:0] select_ln346_186_fu_17709_p3;
wire   [20:0] select_ln346_188_fu_17731_p3;
wire   [20:0] select_ln346_189_fu_17738_p3;
wire   [0:0] tmp_437_fu_17744_p3;
wire   [0:0] tmp_438_fu_17752_p3;
wire   [0:0] xor_ln895_158_fu_17760_p2;
wire   [0:0] and_ln895_114_fu_17766_p2;
wire   [0:0] xor_ln346_24_fu_17780_p2;
wire   [20:0] select_ln346_190_fu_17772_p3;
wire   [20:0] select_ln346_191_fu_17786_p3;
wire   [0:0] tmp_439_fu_17794_p3;
wire   [0:0] tmp_440_fu_17802_p3;
wire   [0:0] xor_ln895_159_fu_17810_p2;
wire   [0:0] and_ln895_115_fu_17816_p2;
wire   [0:0] xor_ln346_25_fu_17830_p2;
wire   [20:0] select_ln346_192_fu_17822_p3;
wire   [20:0] select_ln346_194_fu_17848_p3;
wire  signed [20:0] sext_ln856_5_fu_17845_p1;
wire   [20:0] select_ln346_195_fu_17855_p3;
wire   [0:0] tmp_447_fu_17862_p3;
wire   [0:0] tmp_448_fu_17870_p3;
wire   [0:0] xor_ln895_162_fu_17878_p2;
wire   [0:0] and_ln895_117_fu_17884_p2;
wire   [0:0] xor_ln346_26_fu_17898_p2;
wire   [20:0] select_ln346_196_fu_17890_p3;
wire   [20:0] select_ln346_197_fu_17904_p3;
wire   [0:0] tmp_449_fu_17912_p3;
wire   [0:0] tmp_450_fu_17920_p3;
wire   [0:0] xor_ln895_163_fu_17928_p2;
wire   [0:0] and_ln895_118_fu_17934_p2;
wire   [0:0] xor_ln346_27_fu_17948_p2;
wire   [20:0] select_ln346_198_fu_17940_p3;
wire   [0:0] and_ln378_54_fu_17963_p2;
wire   [0:0] and_ln891_54_fu_17967_p2;
wire   [0:0] xor_ln896_182_fu_17972_p2;
wire   [0:0] and_ln896_54_fu_17977_p2;
wire   [0:0] or_ln346_54_fu_17989_p2;
wire   [20:0] select_ln346_202_fu_17982_p3;
wire   [20:0] select_ln346_203_fu_17994_p3;
wire   [0:0] tmp_463_fu_18001_p3;
wire   [0:0] tmp_464_fu_18009_p3;
wire   [0:0] xor_ln895_168_fu_18017_p2;
wire   [0:0] and_ln895_121_fu_18023_p2;
wire   [0:0] xor_ln346_28_fu_18037_p2;
wire   [20:0] select_ln346_204_fu_18029_p3;
wire   [0:0] and_ln378_56_fu_18051_p2;
wire   [0:0] and_ln891_56_fu_18055_p2;
wire   [0:0] xor_ln896_184_fu_18060_p2;
wire   [0:0] and_ln896_56_fu_18065_p2;
wire   [0:0] or_ln346_56_fu_18077_p2;
wire   [20:0] select_ln346_208_fu_18070_p3;
wire   [20:0] select_ln346_209_fu_18082_p3;
wire   [0:0] tmp_477_fu_18089_p3;
wire   [0:0] tmp_478_fu_18097_p3;
wire   [0:0] xor_ln895_173_fu_18105_p2;
wire   [0:0] and_ln895_124_fu_18111_p2;
wire   [0:0] xor_ln346_29_fu_18125_p2;
wire   [20:0] select_ln346_210_fu_18117_p3;
wire  signed [34:0] shl_ln838_41_fu_18139_p3;
wire  signed [35:0] sext_ln813_119_fu_18146_p1;
wire  signed [35:0] sext_ln1347_59_fu_18150_p1;
wire   [35:0] add_ln1347_60_fu_18153_p2;
(* use_dsp48 = "no" *) wire   [34:0] add_ln810_36_fu_18159_p2;
wire   [20:0] zext_ln377_59_fu_18190_p1;
wire   [20:0] trunc_ln818_58_fu_18172_p4;
wire   [20:0] add_ln377_59_fu_18193_p2;
wire   [0:0] tmp_494_fu_18199_p3;
wire   [0:0] tmp_492_fu_18182_p3;
wire   [0:0] xor_ln896_148_fu_18207_p2;
wire   [0:0] xor_ln888_118_fu_18227_p2;
wire   [0:0] tmp_495_fu_18219_p3;
wire   [0:0] or_ln888_59_fu_18233_p2;
wire   [0:0] tmp_496_fu_18245_p3;
wire   [0:0] xor_ln890_59_fu_18253_p2;
wire   [0:0] or_ln890_59_fu_18259_p2;
wire   [0:0] and_ln378_59_fu_18213_p2;
wire   [0:0] xor_ln888_119_fu_18239_p2;
wire   [0:0] xor_ln895_178_fu_18277_p2;
wire   [0:0] tmp_491_fu_18164_p3;
wire   [0:0] or_ln895_59_fu_18283_p2;
wire   [0:0] xor_ln895_179_fu_18289_p2;
wire   [0:0] and_ln890_59_fu_18265_p2;
wire   [0:0] xor_ln896_149_fu_18301_p2;
wire   [0:0] and_ln891_59_fu_18271_p2;
wire   [0:0] or_ln896_59_fu_18307_p2;
wire   [0:0] xor_ln896_187_fu_18313_p2;
wire   [0:0] and_ln895_127_fu_18295_p2;
wire   [0:0] and_ln896_59_fu_18319_p2;
wire   [0:0] or_ln346_59_fu_18333_p2;
wire   [20:0] select_ln346_216_fu_18325_p3;
wire  signed [34:0] shl_ln838_43_fu_18347_p3;
wire  signed [35:0] sext_ln813_121_fu_18354_p1;
wire  signed [35:0] sext_ln1347_62_fu_18358_p1;
wire  signed [34:0] sext_ln1347_63_fu_18361_p1;
wire   [35:0] add_ln1347_62_fu_18364_p2;
wire   [34:0] add_ln810_38_fu_18370_p2;
wire   [20:0] zext_ln377_62_fu_18402_p1;
wire   [20:0] trunc_ln818_61_fu_18384_p4;
wire   [20:0] add_ln377_62_fu_18405_p2;
wire   [0:0] tmp_512_fu_18411_p3;
wire   [0:0] tmp_510_fu_18394_p3;
wire   [0:0] xor_ln896_154_fu_18419_p2;
wire   [0:0] xor_ln888_124_fu_18439_p2;
wire   [0:0] tmp_513_fu_18431_p3;
wire   [0:0] or_ln888_62_fu_18445_p2;
wire   [0:0] tmp_514_fu_18457_p3;
wire   [0:0] xor_ln890_62_fu_18465_p2;
wire   [0:0] or_ln890_62_fu_18471_p2;
wire   [0:0] and_ln378_62_fu_18425_p2;
wire   [0:0] xor_ln888_125_fu_18451_p2;
wire   [0:0] xor_ln895_184_fu_18489_p2;
wire   [0:0] tmp_509_fu_18376_p3;
wire   [0:0] or_ln895_62_fu_18495_p2;
wire   [0:0] xor_ln895_185_fu_18501_p2;
wire   [0:0] and_ln890_62_fu_18477_p2;
wire   [0:0] xor_ln896_155_fu_18513_p2;
wire   [0:0] and_ln891_62_fu_18483_p2;
wire   [0:0] or_ln896_62_fu_18519_p2;
wire   [0:0] xor_ln896_190_fu_18525_p2;
wire   [0:0] and_ln895_130_fu_18507_p2;
wire   [0:0] and_ln896_62_fu_18531_p2;
wire   [0:0] or_ln346_62_fu_18545_p2;
wire   [20:0] select_ln346_222_fu_18537_p3;
wire  signed [20:0] sext_ln813_123_fu_18563_p0;
wire  signed [21:0] sext_ln813_123_fu_18563_p1;
wire  signed [21:0] sext_ln813_122_fu_18559_p1;
wire   [21:0] add_ln1347_63_fu_18567_p2;
wire  signed [20:0] add_ln813_18_fu_18581_p0;
wire   [20:0] add_ln813_18_fu_18581_p2;
wire   [0:0] tmp_544_fu_18573_p3;
wire   [0:0] tmp_545_fu_18587_p3;
wire   [0:0] xor_ln895_198_fu_18595_p2;
wire   [0:0] and_ln895_143_fu_18601_p2;
wire   [0:0] xor_ln302_24_fu_18607_p2;
wire   [20:0] select_ln346_248_fu_18613_p3;
wire  signed [20:0] sext_ln813_125_fu_18634_p0;
wire  signed [21:0] sext_ln813_125_fu_18634_p1;
wire  signed [21:0] sext_ln813_124_fu_18630_p1;
wire   [21:0] add_ln1347_64_fu_18638_p2;
wire  signed [20:0] add_ln813_19_fu_18652_p0;
wire   [20:0] add_ln813_19_fu_18652_p2;
wire   [0:0] tmp_546_fu_18644_p3;
wire   [0:0] tmp_547_fu_18658_p3;
wire   [0:0] xor_ln895_199_fu_18666_p2;
wire   [0:0] and_ln895_144_fu_18672_p2;
wire   [0:0] xor_ln302_25_fu_18678_p2;
wire   [20:0] select_ln346_249_fu_18684_p3;
wire   [0:0] grp_fu_1188_p2;
wire   [19:0] trunc_ln1649_fu_18701_p1;
wire   [19:0] select_ln49_fu_18705_p3;
wire   [0:0] grp_fu_1194_p2;
wire   [19:0] trunc_ln1649_1_fu_18718_p1;
wire   [19:0] select_ln49_1_fu_18722_p3;
wire  signed [20:0] sext_ln813_127_fu_18739_p0;
wire  signed [21:0] sext_ln813_127_fu_18739_p1;
wire  signed [21:0] sext_ln813_126_fu_18735_p1;
wire   [21:0] add_ln1347_65_fu_18743_p2;
wire  signed [20:0] add_ln813_20_fu_18757_p0;
wire   [20:0] add_ln813_20_fu_18757_p2;
wire   [0:0] tmp_548_fu_18749_p3;
wire   [0:0] tmp_549_fu_18763_p3;
wire   [0:0] xor_ln895_200_fu_18771_p2;
wire   [0:0] and_ln895_145_fu_18777_p2;
wire   [0:0] xor_ln302_26_fu_18783_p2;
wire   [20:0] select_ln346_250_fu_18789_p3;
wire  signed [20:0] sext_ln813_129_fu_18810_p0;
wire  signed [21:0] sext_ln813_129_fu_18810_p1;
wire  signed [21:0] sext_ln813_128_fu_18806_p1;
wire   [21:0] add_ln1347_66_fu_18814_p2;
wire  signed [20:0] add_ln813_21_fu_18828_p0;
wire   [20:0] add_ln813_21_fu_18828_p2;
wire   [0:0] tmp_550_fu_18820_p3;
wire   [0:0] tmp_551_fu_18834_p3;
wire   [0:0] xor_ln895_201_fu_18842_p2;
wire   [0:0] and_ln895_146_fu_18848_p2;
wire   [0:0] xor_ln302_27_fu_18854_p2;
wire   [20:0] select_ln346_251_fu_18860_p3;
wire   [19:0] trunc_ln1649_2_fu_18877_p1;
wire   [19:0] select_ln49_2_fu_18881_p3;
wire   [19:0] trunc_ln1649_3_fu_18894_p1;
wire   [19:0] select_ln49_3_fu_18898_p3;
wire  signed [20:0] sext_ln813_131_fu_18915_p0;
wire  signed [21:0] sext_ln813_131_fu_18915_p1;
wire  signed [21:0] sext_ln813_130_fu_18911_p1;
wire   [21:0] add_ln1347_67_fu_18919_p2;
wire  signed [20:0] add_ln813_22_fu_18933_p0;
wire   [20:0] add_ln813_22_fu_18933_p2;
wire   [0:0] tmp_552_fu_18925_p3;
wire   [0:0] tmp_553_fu_18939_p3;
wire   [0:0] xor_ln895_202_fu_18947_p2;
wire   [0:0] and_ln895_147_fu_18953_p2;
wire   [0:0] xor_ln302_28_fu_18959_p2;
wire   [20:0] select_ln346_252_fu_18965_p3;
wire  signed [20:0] sext_ln813_133_fu_18986_p0;
wire  signed [21:0] sext_ln813_133_fu_18986_p1;
wire  signed [21:0] sext_ln813_132_fu_18982_p1;
wire   [21:0] add_ln1347_68_fu_18990_p2;
wire  signed [20:0] add_ln813_23_fu_19004_p0;
wire   [20:0] add_ln813_23_fu_19004_p2;
wire   [0:0] tmp_554_fu_18996_p3;
wire   [0:0] tmp_555_fu_19010_p3;
wire   [0:0] xor_ln895_203_fu_19018_p2;
wire   [0:0] and_ln895_148_fu_19024_p2;
wire   [0:0] xor_ln302_29_fu_19030_p2;
wire   [20:0] select_ln346_253_fu_19036_p3;
wire   [19:0] trunc_ln1649_4_fu_19053_p1;
wire   [19:0] select_ln49_4_fu_19057_p3;
wire   [19:0] trunc_ln1649_5_fu_19070_p1;
wire   [19:0] select_ln49_5_fu_19074_p3;
wire  signed [20:0] sext_ln813_135_fu_19091_p0;
wire  signed [21:0] sext_ln813_135_fu_19091_p1;
wire  signed [21:0] sext_ln813_134_fu_19087_p1;
wire   [21:0] add_ln1347_69_fu_19095_p2;
wire  signed [20:0] add_ln813_24_fu_19109_p0;
wire   [20:0] add_ln813_24_fu_19109_p2;
wire   [0:0] tmp_556_fu_19101_p3;
wire   [0:0] tmp_557_fu_19115_p3;
wire   [0:0] xor_ln895_204_fu_19123_p2;
wire   [0:0] and_ln895_149_fu_19129_p2;
wire   [0:0] xor_ln302_30_fu_19135_p2;
wire   [20:0] select_ln346_254_fu_19141_p3;
wire  signed [20:0] sext_ln813_137_fu_19162_p0;
wire  signed [21:0] sext_ln813_137_fu_19162_p1;
wire  signed [21:0] sext_ln813_136_fu_19158_p1;
wire   [21:0] add_ln1347_70_fu_19166_p2;
wire  signed [20:0] add_ln813_25_fu_19180_p0;
wire   [20:0] add_ln813_25_fu_19180_p2;
wire   [0:0] tmp_558_fu_19172_p3;
wire   [0:0] tmp_559_fu_19186_p3;
wire   [0:0] xor_ln895_205_fu_19194_p2;
wire   [0:0] and_ln895_150_fu_19200_p2;
wire   [0:0] xor_ln302_31_fu_19206_p2;
wire   [20:0] select_ln346_255_fu_19212_p3;
wire   [19:0] trunc_ln1649_6_fu_19229_p1;
wire   [19:0] select_ln49_6_fu_19233_p3;
wire   [19:0] trunc_ln1649_7_fu_19246_p1;
wire   [19:0] select_ln49_7_fu_19250_p3;
wire  signed [20:0] sext_ln813_139_fu_19267_p0;
wire  signed [21:0] sext_ln813_139_fu_19267_p1;
wire  signed [21:0] sext_ln813_138_fu_19263_p1;
wire   [21:0] add_ln1347_71_fu_19271_p2;
wire  signed [20:0] add_ln813_26_fu_19285_p0;
wire   [20:0] add_ln813_26_fu_19285_p2;
wire   [0:0] tmp_560_fu_19277_p3;
wire   [0:0] tmp_561_fu_19291_p3;
wire   [0:0] xor_ln895_206_fu_19299_p2;
wire   [0:0] and_ln895_151_fu_19305_p2;
wire   [0:0] xor_ln302_32_fu_19311_p2;
wire   [20:0] select_ln346_256_fu_19317_p3;
wire  signed [20:0] sext_ln813_141_fu_19338_p0;
wire  signed [21:0] sext_ln813_141_fu_19338_p1;
wire  signed [21:0] sext_ln813_140_fu_19334_p1;
wire   [21:0] add_ln1347_72_fu_19342_p2;
wire  signed [20:0] add_ln813_27_fu_19356_p0;
wire   [20:0] add_ln813_27_fu_19356_p2;
wire   [0:0] tmp_562_fu_19348_p3;
wire   [0:0] tmp_563_fu_19362_p3;
wire   [0:0] xor_ln895_207_fu_19370_p2;
wire   [0:0] and_ln895_152_fu_19376_p2;
wire   [0:0] xor_ln302_33_fu_19382_p2;
wire   [20:0] select_ln346_257_fu_19388_p3;
wire   [19:0] trunc_ln1649_8_fu_19405_p1;
wire   [19:0] select_ln49_8_fu_19409_p3;
wire   [19:0] trunc_ln1649_9_fu_19422_p1;
wire   [19:0] select_ln49_9_fu_19426_p3;
wire  signed [20:0] sext_ln813_143_fu_19443_p0;
wire  signed [21:0] sext_ln813_143_fu_19443_p1;
wire  signed [21:0] sext_ln813_142_fu_19439_p1;
wire   [21:0] add_ln1347_73_fu_19447_p2;
wire  signed [20:0] add_ln813_28_fu_19461_p0;
wire   [20:0] add_ln813_28_fu_19461_p2;
wire   [0:0] tmp_564_fu_19453_p3;
wire   [0:0] tmp_565_fu_19467_p3;
wire   [0:0] xor_ln895_208_fu_19475_p2;
wire   [0:0] and_ln895_153_fu_19481_p2;
wire   [0:0] xor_ln302_34_fu_19487_p2;
wire   [20:0] select_ln346_258_fu_19493_p3;
wire  signed [20:0] sext_ln813_145_fu_19514_p0;
wire  signed [21:0] sext_ln813_145_fu_19514_p1;
wire  signed [21:0] sext_ln813_144_fu_19510_p1;
wire   [21:0] add_ln1347_74_fu_19518_p2;
wire  signed [20:0] add_ln813_29_fu_19532_p0;
wire   [20:0] add_ln813_29_fu_19532_p2;
wire   [0:0] tmp_566_fu_19524_p3;
wire   [0:0] tmp_567_fu_19538_p3;
wire   [0:0] xor_ln895_209_fu_19546_p2;
wire   [0:0] and_ln895_154_fu_19552_p2;
wire   [0:0] xor_ln302_35_fu_19558_p2;
wire   [20:0] select_ln346_259_fu_19564_p3;
wire   [19:0] trunc_ln1649_10_fu_19581_p1;
wire   [19:0] select_ln49_10_fu_19585_p3;
wire   [19:0] trunc_ln1649_11_fu_19598_p1;
wire   [19:0] select_ln49_11_fu_19602_p3;
wire  signed [20:0] sext_ln813_147_fu_19619_p0;
wire  signed [21:0] sext_ln813_147_fu_19619_p1;
wire  signed [21:0] sext_ln813_146_fu_19615_p1;
wire   [21:0] add_ln1347_75_fu_19623_p2;
wire  signed [20:0] add_ln813_30_fu_19637_p0;
wire   [20:0] add_ln813_30_fu_19637_p2;
wire   [0:0] tmp_568_fu_19629_p3;
wire   [0:0] tmp_569_fu_19643_p3;
wire   [0:0] xor_ln895_210_fu_19651_p2;
wire   [0:0] and_ln895_155_fu_19657_p2;
wire   [0:0] xor_ln302_36_fu_19663_p2;
wire   [20:0] select_ln346_260_fu_19669_p3;
wire  signed [20:0] sext_ln813_149_fu_19690_p0;
wire  signed [21:0] sext_ln813_149_fu_19690_p1;
wire  signed [21:0] sext_ln813_148_fu_19686_p1;
wire   [21:0] add_ln1347_76_fu_19694_p2;
wire  signed [20:0] add_ln813_31_fu_19708_p0;
wire   [20:0] add_ln813_31_fu_19708_p2;
wire   [0:0] tmp_570_fu_19700_p3;
wire   [0:0] tmp_571_fu_19714_p3;
wire   [0:0] xor_ln895_211_fu_19722_p2;
wire   [0:0] and_ln895_156_fu_19728_p2;
wire   [0:0] xor_ln302_37_fu_19734_p2;
wire   [20:0] select_ln346_261_fu_19740_p3;
wire   [19:0] trunc_ln1649_12_fu_19757_p1;
wire   [19:0] select_ln49_12_fu_19761_p3;
wire   [19:0] trunc_ln1649_13_fu_19774_p1;
wire   [19:0] select_ln49_13_fu_19778_p3;
wire  signed [20:0] sext_ln813_151_fu_19795_p0;
wire  signed [21:0] sext_ln813_151_fu_19795_p1;
wire  signed [21:0] sext_ln813_150_fu_19791_p1;
wire   [21:0] add_ln1347_77_fu_19799_p2;
wire  signed [20:0] add_ln813_32_fu_19813_p0;
wire   [20:0] add_ln813_32_fu_19813_p2;
wire   [0:0] tmp_572_fu_19805_p3;
wire   [0:0] tmp_573_fu_19819_p3;
wire   [0:0] xor_ln895_212_fu_19827_p2;
wire   [0:0] and_ln895_157_fu_19833_p2;
wire   [0:0] xor_ln302_38_fu_19839_p2;
wire   [20:0] select_ln346_262_fu_19845_p3;
wire  signed [20:0] sext_ln813_153_fu_19866_p0;
wire  signed [21:0] sext_ln813_153_fu_19866_p1;
wire  signed [21:0] sext_ln813_152_fu_19862_p1;
wire   [21:0] add_ln1347_78_fu_19870_p2;
wire  signed [20:0] add_ln813_33_fu_19884_p0;
wire   [20:0] add_ln813_33_fu_19884_p2;
wire   [0:0] tmp_574_fu_19876_p3;
wire   [0:0] tmp_575_fu_19890_p3;
wire   [0:0] xor_ln895_213_fu_19898_p2;
wire   [0:0] and_ln895_158_fu_19904_p2;
wire   [0:0] xor_ln302_39_fu_19910_p2;
wire   [20:0] select_ln346_263_fu_19916_p3;
wire   [19:0] trunc_ln1649_14_fu_19933_p1;
wire   [19:0] select_ln49_14_fu_19937_p3;
wire   [19:0] trunc_ln1649_15_fu_19950_p1;
wire   [19:0] select_ln49_15_fu_19954_p3;
wire  signed [20:0] sext_ln813_155_fu_19971_p0;
wire  signed [21:0] sext_ln813_155_fu_19971_p1;
wire  signed [21:0] sext_ln813_154_fu_19967_p1;
wire   [21:0] add_ln1347_79_fu_19975_p2;
wire  signed [20:0] add_ln813_34_fu_19989_p0;
wire   [20:0] add_ln813_34_fu_19989_p2;
wire   [0:0] tmp_576_fu_19981_p3;
wire   [0:0] tmp_577_fu_19995_p3;
wire   [0:0] xor_ln895_214_fu_20003_p2;
wire   [0:0] and_ln895_159_fu_20009_p2;
wire   [0:0] xor_ln302_40_fu_20015_p2;
wire   [20:0] select_ln346_264_fu_20021_p3;
wire  signed [20:0] sext_ln813_157_fu_20042_p0;
wire  signed [21:0] sext_ln813_157_fu_20042_p1;
wire  signed [21:0] sext_ln813_156_fu_20038_p1;
wire   [21:0] add_ln1347_80_fu_20046_p2;
wire  signed [20:0] add_ln813_35_fu_20060_p0;
wire   [20:0] add_ln813_35_fu_20060_p2;
wire   [0:0] tmp_578_fu_20052_p3;
wire   [0:0] tmp_579_fu_20066_p3;
wire   [0:0] xor_ln895_215_fu_20074_p2;
wire   [0:0] and_ln895_160_fu_20080_p2;
wire   [0:0] xor_ln302_41_fu_20086_p2;
wire   [20:0] select_ln346_265_fu_20092_p3;
wire   [19:0] trunc_ln1649_16_fu_20109_p1;
wire   [19:0] select_ln49_16_fu_20113_p3;
wire   [19:0] trunc_ln1649_17_fu_20126_p1;
wire   [19:0] select_ln49_17_fu_20130_p3;
wire  signed [20:0] sext_ln813_158_fu_20143_p0;
wire  signed [21:0] sext_ln813_159_fu_20147_p1;
wire  signed [21:0] sext_ln813_158_fu_20143_p1;
wire   [21:0] add_ln1347_81_fu_20150_p2;
wire  signed [20:0] add_ln813_36_fu_20164_p1;
wire   [20:0] add_ln813_36_fu_20164_p2;
wire   [0:0] tmp_580_fu_20156_p3;
wire   [0:0] tmp_581_fu_20169_p3;
wire   [0:0] xor_ln895_216_fu_20177_p2;
wire   [0:0] and_ln895_161_fu_20183_p2;
wire   [0:0] xor_ln302_42_fu_20189_p2;
wire   [20:0] select_ln346_266_fu_20195_p3;
wire  signed [20:0] sext_ln813_160_fu_20212_p0;
wire  signed [21:0] sext_ln813_161_fu_20216_p1;
wire  signed [21:0] sext_ln813_160_fu_20212_p1;
wire   [21:0] add_ln1347_82_fu_20219_p2;
wire  signed [20:0] add_ln813_37_fu_20233_p1;
wire   [20:0] add_ln813_37_fu_20233_p2;
wire   [0:0] tmp_582_fu_20225_p3;
wire   [0:0] tmp_583_fu_20238_p3;
wire   [0:0] xor_ln895_217_fu_20246_p2;
wire   [0:0] and_ln895_162_fu_20252_p2;
wire   [0:0] xor_ln302_43_fu_20258_p2;
wire   [20:0] select_ln346_267_fu_20264_p3;
wire  signed [20:0] sext_ln813_162_fu_20281_p0;
wire  signed [21:0] sext_ln813_163_fu_20285_p1;
wire  signed [21:0] sext_ln813_162_fu_20281_p1;
wire   [21:0] add_ln1347_83_fu_20288_p2;
wire  signed [20:0] add_ln813_38_fu_20302_p1;
wire   [20:0] add_ln813_38_fu_20302_p2;
wire   [0:0] tmp_584_fu_20294_p3;
wire   [0:0] tmp_585_fu_20307_p3;
wire   [0:0] xor_ln895_218_fu_20315_p2;
wire   [0:0] and_ln895_163_fu_20321_p2;
wire   [0:0] xor_ln302_44_fu_20327_p2;
wire   [20:0] select_ln346_268_fu_20333_p3;
wire  signed [20:0] sext_ln813_164_fu_20350_p0;
wire  signed [21:0] sext_ln813_165_fu_20354_p1;
wire  signed [21:0] sext_ln813_164_fu_20350_p1;
wire   [21:0] add_ln1347_84_fu_20357_p2;
wire  signed [20:0] add_ln813_39_fu_20371_p1;
wire   [20:0] add_ln813_39_fu_20371_p2;
wire   [0:0] tmp_586_fu_20363_p3;
wire   [0:0] tmp_587_fu_20376_p3;
wire   [0:0] xor_ln895_219_fu_20384_p2;
wire   [0:0] and_ln895_164_fu_20390_p2;
wire   [0:0] xor_ln302_45_fu_20396_p2;
wire   [20:0] select_ln346_269_fu_20402_p3;
wire  signed [20:0] sext_ln813_166_fu_20419_p0;
wire  signed [21:0] sext_ln813_167_fu_20423_p1;
wire  signed [21:0] sext_ln813_166_fu_20419_p1;
wire   [21:0] add_ln1347_85_fu_20426_p2;
wire  signed [20:0] add_ln813_40_fu_20440_p1;
wire   [20:0] add_ln813_40_fu_20440_p2;
wire   [0:0] tmp_588_fu_20432_p3;
wire   [0:0] tmp_589_fu_20445_p3;
wire   [0:0] xor_ln895_220_fu_20453_p2;
wire   [0:0] and_ln895_165_fu_20459_p2;
wire   [0:0] xor_ln302_46_fu_20465_p2;
wire   [20:0] select_ln346_270_fu_20471_p3;
wire  signed [20:0] sext_ln813_168_fu_20488_p0;
wire  signed [21:0] sext_ln813_169_fu_20492_p1;
wire  signed [21:0] sext_ln813_168_fu_20488_p1;
wire   [21:0] add_ln1347_86_fu_20495_p2;
wire  signed [20:0] add_ln813_41_fu_20509_p1;
wire   [20:0] add_ln813_41_fu_20509_p2;
wire   [0:0] tmp_590_fu_20501_p3;
wire   [0:0] tmp_591_fu_20514_p3;
wire   [0:0] xor_ln895_221_fu_20522_p2;
wire   [0:0] and_ln895_166_fu_20528_p2;
wire   [0:0] xor_ln302_47_fu_20534_p2;
wire   [20:0] select_ln346_271_fu_20540_p3;
wire  signed [20:0] sext_ln813_170_fu_20557_p0;
wire  signed [21:0] sext_ln813_171_fu_20561_p1;
wire  signed [21:0] sext_ln813_170_fu_20557_p1;
wire   [21:0] add_ln1347_87_fu_20564_p2;
wire  signed [20:0] add_ln813_42_fu_20578_p1;
wire   [20:0] add_ln813_42_fu_20578_p2;
wire   [0:0] tmp_592_fu_20570_p3;
wire   [0:0] tmp_593_fu_20583_p3;
wire   [0:0] xor_ln895_222_fu_20591_p2;
wire   [0:0] and_ln895_167_fu_20597_p2;
wire   [0:0] xor_ln302_48_fu_20603_p2;
wire   [20:0] select_ln346_272_fu_20609_p3;
wire  signed [20:0] sext_ln813_172_fu_20626_p0;
wire  signed [21:0] sext_ln813_173_fu_20630_p1;
wire  signed [21:0] sext_ln813_172_fu_20626_p1;
wire   [21:0] add_ln1347_88_fu_20633_p2;
wire  signed [20:0] add_ln813_43_fu_20647_p1;
wire   [20:0] add_ln813_43_fu_20647_p2;
wire   [0:0] tmp_594_fu_20639_p3;
wire   [0:0] tmp_595_fu_20652_p3;
wire   [0:0] xor_ln895_223_fu_20660_p2;
wire   [0:0] and_ln895_168_fu_20666_p2;
wire   [0:0] xor_ln302_49_fu_20672_p2;
wire   [20:0] select_ln346_273_fu_20678_p3;
wire  signed [20:0] sext_ln813_174_fu_20695_p0;
wire  signed [21:0] sext_ln813_175_fu_20699_p1;
wire  signed [21:0] sext_ln813_174_fu_20695_p1;
wire   [21:0] add_ln1347_89_fu_20702_p2;
wire  signed [20:0] add_ln813_44_fu_20716_p1;
wire   [20:0] add_ln813_44_fu_20716_p2;
wire   [0:0] tmp_596_fu_20708_p3;
wire   [0:0] tmp_597_fu_20721_p3;
wire   [0:0] xor_ln895_224_fu_20729_p2;
wire   [0:0] and_ln895_169_fu_20735_p2;
wire   [0:0] xor_ln302_50_fu_20741_p2;
wire   [20:0] select_ln346_274_fu_20747_p3;
wire  signed [20:0] sext_ln813_176_fu_20764_p0;
wire  signed [21:0] sext_ln813_177_fu_20768_p1;
wire  signed [21:0] sext_ln813_176_fu_20764_p1;
wire   [21:0] add_ln1347_90_fu_20771_p2;
wire  signed [20:0] add_ln813_45_fu_20785_p1;
wire   [20:0] add_ln813_45_fu_20785_p2;
wire   [0:0] tmp_598_fu_20777_p3;
wire   [0:0] tmp_599_fu_20790_p3;
wire   [0:0] xor_ln895_225_fu_20798_p2;
wire   [0:0] and_ln895_170_fu_20804_p2;
wire   [0:0] xor_ln302_51_fu_20810_p2;
wire   [20:0] select_ln346_275_fu_20816_p3;
wire  signed [20:0] sext_ln813_178_fu_20833_p0;
wire  signed [21:0] sext_ln813_179_fu_20837_p1;
wire  signed [21:0] sext_ln813_178_fu_20833_p1;
wire   [21:0] add_ln1347_91_fu_20840_p2;
wire  signed [20:0] add_ln813_46_fu_20854_p1;
wire   [20:0] add_ln813_46_fu_20854_p2;
wire   [0:0] tmp_600_fu_20846_p3;
wire   [0:0] tmp_601_fu_20859_p3;
wire   [0:0] xor_ln895_226_fu_20867_p2;
wire   [0:0] and_ln895_171_fu_20873_p2;
wire   [0:0] xor_ln302_52_fu_20879_p2;
wire   [20:0] select_ln346_276_fu_20885_p3;
wire  signed [20:0] sext_ln813_180_fu_20902_p0;
wire  signed [21:0] sext_ln813_181_fu_20906_p1;
wire  signed [21:0] sext_ln813_180_fu_20902_p1;
wire   [21:0] add_ln1347_92_fu_20909_p2;
wire  signed [20:0] add_ln813_47_fu_20923_p1;
wire   [20:0] add_ln813_47_fu_20923_p2;
wire   [0:0] tmp_602_fu_20915_p3;
wire   [0:0] tmp_603_fu_20928_p3;
wire   [0:0] xor_ln895_227_fu_20936_p2;
wire   [0:0] and_ln895_172_fu_20942_p2;
wire   [0:0] xor_ln302_53_fu_20948_p2;
wire   [20:0] select_ln346_277_fu_20954_p3;
wire  signed [20:0] sext_ln813_182_fu_20971_p0;
wire  signed [21:0] sext_ln813_183_fu_20975_p1;
wire  signed [21:0] sext_ln813_182_fu_20971_p1;
wire   [21:0] add_ln1347_93_fu_20978_p2;
wire  signed [20:0] add_ln813_48_fu_20992_p1;
wire   [20:0] add_ln813_48_fu_20992_p2;
wire   [0:0] tmp_604_fu_20984_p3;
wire   [0:0] tmp_605_fu_20997_p3;
wire   [0:0] xor_ln895_228_fu_21005_p2;
wire   [0:0] and_ln895_173_fu_21011_p2;
wire   [0:0] xor_ln302_54_fu_21017_p2;
wire   [20:0] select_ln346_278_fu_21023_p3;
wire  signed [20:0] sext_ln813_184_fu_21040_p0;
wire  signed [21:0] sext_ln813_185_fu_21044_p1;
wire  signed [21:0] sext_ln813_184_fu_21040_p1;
wire   [21:0] add_ln1347_94_fu_21047_p2;
wire  signed [20:0] add_ln813_49_fu_21061_p1;
wire   [20:0] add_ln813_49_fu_21061_p2;
wire   [0:0] tmp_606_fu_21053_p3;
wire   [0:0] tmp_607_fu_21066_p3;
wire   [0:0] xor_ln895_229_fu_21074_p2;
wire   [0:0] and_ln895_174_fu_21080_p2;
wire   [0:0] xor_ln302_55_fu_21086_p2;
wire   [20:0] select_ln346_279_fu_21092_p3;
wire  signed [20:0] sext_ln813_186_fu_21109_p0;
wire  signed [21:0] sext_ln813_187_fu_21113_p1;
wire  signed [21:0] sext_ln813_186_fu_21109_p1;
wire   [21:0] add_ln1347_95_fu_21116_p2;
wire  signed [20:0] add_ln813_50_fu_21130_p1;
wire   [20:0] add_ln813_50_fu_21130_p2;
wire   [0:0] tmp_608_fu_21122_p3;
wire   [0:0] tmp_609_fu_21135_p3;
wire   [0:0] xor_ln895_230_fu_21143_p2;
wire   [0:0] and_ln895_175_fu_21149_p2;
wire   [0:0] xor_ln302_56_fu_21155_p2;
wire   [20:0] select_ln346_280_fu_21161_p3;
wire  signed [20:0] sext_ln813_188_fu_21178_p0;
wire  signed [21:0] sext_ln813_189_fu_21182_p1;
wire  signed [21:0] sext_ln813_188_fu_21178_p1;
wire   [21:0] add_ln1347_96_fu_21185_p2;
wire  signed [20:0] add_ln813_51_fu_21199_p1;
wire   [20:0] add_ln813_51_fu_21199_p2;
wire   [0:0] tmp_610_fu_21191_p3;
wire   [0:0] tmp_611_fu_21204_p3;
wire   [0:0] xor_ln895_231_fu_21212_p2;
wire   [0:0] and_ln895_176_fu_21218_p2;
wire   [0:0] xor_ln302_57_fu_21224_p2;
wire   [20:0] select_ln346_281_fu_21230_p3;
wire  signed [20:0] sext_ln813_190_fu_21247_p0;
wire  signed [21:0] sext_ln813_191_fu_21251_p1;
wire  signed [21:0] sext_ln813_190_fu_21247_p1;
wire   [21:0] add_ln1347_97_fu_21254_p2;
wire  signed [20:0] add_ln813_52_fu_21268_p1;
wire   [20:0] add_ln813_52_fu_21268_p2;
wire   [0:0] tmp_612_fu_21260_p3;
wire   [0:0] tmp_613_fu_21273_p3;
wire   [0:0] xor_ln895_232_fu_21281_p2;
wire   [0:0] and_ln895_177_fu_21287_p2;
wire   [0:0] xor_ln302_58_fu_21293_p2;
wire   [20:0] select_ln346_282_fu_21299_p3;
wire  signed [20:0] sext_ln813_192_fu_21316_p0;
wire  signed [21:0] sext_ln813_193_fu_21320_p1;
wire  signed [21:0] sext_ln813_192_fu_21316_p1;
wire   [21:0] add_ln1347_98_fu_21323_p2;
wire  signed [20:0] add_ln813_53_fu_21337_p1;
wire   [20:0] add_ln813_53_fu_21337_p2;
wire   [0:0] tmp_614_fu_21329_p3;
wire   [0:0] tmp_615_fu_21342_p3;
wire   [0:0] xor_ln895_233_fu_21350_p2;
wire   [0:0] and_ln895_178_fu_21356_p2;
wire   [0:0] xor_ln302_59_fu_21362_p2;
wire   [20:0] select_ln346_283_fu_21368_p3;
wire  signed [13:0] grp_fu_21385_p1;
wire  signed [6:0] grp_fu_21397_p1;
wire  signed [20:0] grp_fu_21404_p0;
wire  signed [13:0] grp_fu_21404_p1;
wire  signed [12:0] grp_fu_21411_p1;
wire  signed [20:0] grp_fu_21418_p0;
wire  signed [13:0] grp_fu_21418_p1;
wire  signed [20:0] grp_fu_21430_p0;
wire  signed [13:0] grp_fu_21430_p1;
wire  signed [20:0] grp_fu_21437_p0;
wire  signed [13:0] grp_fu_21437_p1;
wire  signed [8:0] grp_fu_21449_p1;
wire  signed [6:0] grp_fu_21456_p1;
wire  signed [6:0] grp_fu_21465_p1;
wire   [12:0] grp_fu_21474_p1;
wire   [5:0] grp_fu_21481_p1;
wire  signed [20:0] grp_fu_21488_p0;
wire   [12:0] grp_fu_21488_p1;
wire  signed [20:0] grp_fu_21495_p0;
wire   [12:0] grp_fu_21495_p1;
wire   [5:0] grp_fu_21502_p1;
wire   [11:0] grp_fu_21509_p1;
wire   [7:0] grp_fu_21516_p1;
wire  signed [20:0] grp_fu_21523_p0;
wire   [12:0] grp_fu_21523_p1;
wire  signed [20:0] grp_fu_21530_p0;
wire   [12:0] grp_fu_21530_p1;
wire   [5:0] grp_fu_21539_p1;
wire  signed [14:0] grp_fu_21546_p1;
wire  signed [14:0] grp_fu_21553_p1;
wire   [13:0] grp_fu_21560_p1;
wire  signed [14:0] grp_fu_21567_p1;
wire   [13:0] grp_fu_21575_p1;
wire   [13:0] grp_fu_21582_p1;
wire  signed [20:0] grp_fu_21590_p0;
wire  signed [8:0] grp_fu_21590_p1;
wire   [12:0] grp_fu_21597_p1;
wire  signed [9:0] grp_fu_21604_p1;
wire   [11:0] grp_fu_21611_p1;
wire   [11:0] grp_fu_21618_p1;
wire  signed [9:0] grp_fu_21630_p1;
wire  signed [8:0] grp_fu_21642_p1;
wire  signed [20:0] grp_fu_21654_p0;
wire   [12:0] grp_fu_21654_p1;
wire   [5:0] grp_fu_21666_p1;
wire  signed [20:0] grp_fu_21678_p0;
wire   [12:0] grp_fu_21678_p1;
wire  signed [20:0] grp_fu_21690_p0;
wire   [6:0] grp_fu_21690_p1;
wire  signed [20:0] grp_fu_21702_p0;
wire   [11:0] grp_fu_21702_p1;
wire  signed [20:0] grp_fu_21714_p0;
wire   [12:0] grp_fu_21714_p1;
wire  signed [20:0] grp_fu_21721_p0;
wire   [7:0] grp_fu_21721_p1;
wire  signed [20:0] grp_fu_21733_p0;
wire   [6:0] grp_fu_21733_p1;
wire  signed [20:0] grp_fu_21740_p0;
wire  signed [13:0] grp_fu_21740_p1;
wire  signed [20:0] grp_fu_21752_p0;
wire  signed [7:0] grp_fu_21752_p1;
wire  signed [20:0] grp_fu_21764_p0;
wire  signed [12:0] grp_fu_21764_p1;
wire  signed [20:0] grp_fu_21776_p0;
wire  signed [13:0] grp_fu_21776_p1;
wire  signed [20:0] grp_fu_21783_p0;
wire  signed [8:0] grp_fu_21783_p1;
wire  signed [20:0] grp_fu_21795_p0;
wire  signed [7:0] grp_fu_21795_p1;
wire  signed [20:0] grp_fu_21802_p0;
wire   [12:0] grp_fu_21802_p1;
wire  signed [20:0] grp_fu_21810_p0;
wire   [5:0] grp_fu_21810_p1;
wire  signed [20:0] grp_fu_21819_p0;
wire   [12:0] grp_fu_21819_p1;
wire  signed [20:0] grp_fu_21826_p0;
wire   [5:0] grp_fu_21826_p1;
wire  signed [20:0] grp_fu_21833_p0;
wire  signed [13:0] grp_fu_21833_p1;
wire  signed [20:0] grp_fu_21844_p0;
wire  signed [6:0] grp_fu_21844_p1;
wire  signed [20:0] grp_fu_21855_p0;
wire  signed [13:0] grp_fu_21855_p1;
wire  signed [20:0] grp_fu_21863_p0;
wire  signed [6:0] grp_fu_21863_p1;
wire  signed [20:0] grp_fu_21872_p0;
wire  signed [13:0] grp_fu_21872_p1;
wire  signed [20:0] grp_fu_21879_p0;
wire  signed [6:0] grp_fu_21879_p1;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_ST_fsm_state1_blk;
wire    ap_ST_fsm_state2_blk;
wire    ap_ST_fsm_state3_blk;
wire    ap_ST_fsm_state4_blk;
wire    ap_ST_fsm_state5_blk;
wire    ap_ST_fsm_state6_blk;
wire    ap_ST_fsm_state7_blk;
wire    ap_ST_fsm_state8_blk;
wire    ap_ST_fsm_state9_blk;
wire    ap_ST_fsm_state10_blk;
wire    ap_block_state11_pp0_stage10_iter0;
wire    ap_ST_fsm_state11_blk;
wire    ap_ST_fsm_state12_blk;
wire    ap_ST_fsm_state13_blk;
wire    ap_ST_fsm_state14_blk;
wire    ap_ST_fsm_state15_blk;
wire    ap_ST_fsm_state16_blk;
wire    ap_ST_fsm_state17_blk;
wire    ap_ST_fsm_state18_blk;
wire    ap_ST_fsm_state19_blk;
wire    ap_ST_fsm_state20_blk;
wire    ap_ST_fsm_state21_blk;
wire    ap_ST_fsm_state22_blk;
wire    ap_ST_fsm_state23_blk;
wire    ap_ST_fsm_state24_blk;
wire    ap_ST_fsm_state25_blk;
wire    ap_ST_fsm_state26_blk;
wire    ap_ST_fsm_state27_blk;
wire    ap_ST_fsm_state28_blk;
wire    ap_ST_fsm_state29_blk;
wire    ap_ST_fsm_state30_blk;
wire    ap_ST_fsm_state31_blk;
wire    ap_block_state32_pp0_stage31_iter0;
wire    ap_ST_fsm_state32_blk;
wire    ap_ST_fsm_state33_blk;
wire    ap_ST_fsm_state34_blk;
wire    ap_ST_fsm_state35_blk;
wire    ap_ST_fsm_state36_blk;
wire    ap_ST_fsm_state37_blk;
wire    ap_ST_fsm_state38_blk;
wire    ap_ST_fsm_state39_blk;
wire    ap_ST_fsm_state40_blk;
wire    ap_ST_fsm_state41_blk;
wire    ap_ST_fsm_state42_blk;
wire    ap_ST_fsm_state43_blk;
wire    ap_ST_fsm_state44_blk;
wire    ap_ST_fsm_state45_blk;
wire    ap_block_state46_pp0_stage45_iter0;
wire    ap_ST_fsm_state46_blk;
wire    ap_block_state47_pp0_stage46_iter0;
wire    ap_ST_fsm_state47_blk;
wire    ap_block_state48_pp0_stage47_iter0;
wire    ap_ST_fsm_state48_blk;
wire    ap_block_state49_pp0_stage48_iter0;
wire    ap_ST_fsm_state49_blk;
wire    ap_block_state50_pp0_stage49_iter0;
wire    ap_ST_fsm_state50_blk;
wire    ap_block_state51_pp0_stage50_iter0;
wire    ap_ST_fsm_state51_blk;
wire    ap_block_state52_pp0_stage51_iter0;
wire    ap_ST_fsm_state52_blk;
wire    ap_block_state53_pp0_stage52_iter0;
wire    ap_ST_fsm_state53_blk;
wire    ap_block_state54_pp0_stage53_iter0;
wire    ap_ST_fsm_state54_blk;
wire    ap_block_state55_pp0_stage54_iter0;
wire    ap_ST_fsm_state55_blk;
wire    ap_ST_fsm_state56_blk;
wire    ap_ST_fsm_state57_blk;
wire    ap_ST_fsm_state58_blk;
wire    ap_ST_fsm_state59_blk;
wire    ap_ST_fsm_state60_blk;
wire    ap_ST_fsm_state61_blk;
wire    ap_ST_fsm_state62_blk;
wire    ap_ST_fsm_state63_blk;
wire    ap_ST_fsm_state64_blk;
wire    ap_ST_fsm_state65_blk;
wire    ap_ST_fsm_state66_blk;
wire    ap_ST_fsm_state67_blk;
wire    ap_ST_fsm_state68_blk;
wire    ap_ST_fsm_state69_blk;
wire    ap_ST_fsm_state70_blk;
wire    ap_ST_fsm_state71_blk;
wire    ap_ST_fsm_state72_blk;
wire    ap_ST_fsm_state73_blk;
wire    ap_ST_fsm_state74_blk;
wire    ap_ST_fsm_state75_blk;
wire    ap_ST_fsm_state76_blk;
wire    ap_ST_fsm_state77_blk;
wire    ap_ST_fsm_state78_blk;
wire    ap_ST_fsm_state79_blk;
wire    ap_ST_fsm_state80_blk;
wire    ap_ST_fsm_state81_blk;
wire    ap_ST_fsm_state82_blk;
wire    ap_ST_fsm_state83_blk;
wire    ap_ST_fsm_state84_blk;
wire    ap_ST_fsm_state85_blk;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 85'd1;
#0 grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg = 1'b0;
#0 ap_done_reg = 1'b0;
end

mpc_qp_admm_zk_admm_V_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
zk_admm_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(zk_admm_V_address0),
    .ce0(zk_admm_V_ce0),
    .we0(zk_admm_V_we0),
    .d0(zk_admm_V_d0),
    .q0(zk_admm_V_q0),
    .address1(zk_admm_V_address1),
    .ce1(zk_admm_V_ce1),
    .we1(zk_admm_V_we1),
    .d1(zk_admm_V_d1),
    .q1(zk_admm_V_q1)
);

mpc_qp_admm_zk_admm_V_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
uk_admm_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(uk_admm_V_address0),
    .ce0(uk_admm_V_ce0),
    .we0(uk_admm_V_we0),
    .d0(uk_admm_V_d0),
    .q0(uk_admm_V_q0),
    .address1(uk_admm_V_address1),
    .ce1(uk_admm_V_ce1),
    .we1(uk_admm_V_we1),
    .d1(uk_admm_V_d1),
    .q1(uk_admm_V_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
temp_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(temp_address0),
    .ce0(temp_ce0),
    .we0(temp_we0),
    .d0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0),
    .q0(temp_q0),
    .address1(temp_address1),
    .ce1(temp_ce1),
    .we1(temp_we1),
    .d1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1),
    .q1(temp_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
Hxk_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(Hxk_V_address0),
    .ce0(Hxk_V_ce0),
    .we0(Hxk_V_we0),
    .d0(Hxk_V_d0),
    .q0(Hxk_V_q0),
    .address1(Hxk_V_address1),
    .ce1(Hxk_V_ce1),
    .we1(Hxk_V_we1),
    .d1(Hxk_V_d1),
    .q1(Hxk_V_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
temp4_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(temp4_V_address0),
    .ce0(temp4_V_ce0),
    .we0(temp4_V_we0),
    .d0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0),
    .q0(temp4_V_q0),
    .address1(temp4_V_address1),
    .ce1(temp4_V_ce1),
    .we1(temp4_V_we1),
    .d1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1),
    .q1(temp4_V_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
temp5_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(temp5_address0),
    .ce0(temp5_ce0),
    .we0(temp5_we0),
    .d0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0),
    .q0(temp5_q0),
    .address1(temp5_address1),
    .ce1(temp5_ce1),
    .we1(temp5_we1),
    .d1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1),
    .q1(temp5_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
temp6_V_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(temp6_V_address0),
    .ce0(temp6_V_ce0),
    .we0(temp6_V_we0),
    .d0(temp6_V_d0),
    .q0(temp6_V_q0),
    .address1(temp6_V_address1),
    .ce1(temp6_V_ce1),
    .we1(temp6_V_we1),
    .d1(temp6_V_d1),
    .q1(temp6_V_q1)
);

mpc_qp_admm_temp_RAM_AUTO_1R1W #(
    .DataWidth( 21 ),
    .AddressRange( 18 ),
    .AddressWidth( 5 ))
temp7_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(temp7_address0),
    .ce0(temp7_ce0),
    .we0(temp7_we0),
    .d0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0),
    .q0(temp7_q0),
    .address1(temp7_address1),
    .ce1(temp7_ce1),
    .we1(temp7_we1),
    .d1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1),
    .q1(temp7_q1)
);

mpc_vsub_18_ap_fixed_21_7_0_0_0_s grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start),
    .ap_done(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_done),
    .ap_idle(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_idle),
    .ap_ready(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_ready),
    .ap_ce(1'b1),
    .A_address0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0),
    .A_ce0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0),
    .A_q0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0),
    .A_address1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1),
    .A_ce1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1),
    .A_q1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1),
    .B_address0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address0),
    .B_ce0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce0),
    .B_q0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0),
    .B_address1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address1),
    .B_ce1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce1),
    .B_q1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1),
    .R_address0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0),
    .R_ce0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0),
    .R_we0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0),
    .R_d0(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d0),
    .R_address1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1),
    .R_ce1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1),
    .R_we1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1),
    .R_d1(grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_d1)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U42(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_fu_1371_p3),
    .din1(grp_fu_21385_p1),
    .ce(1'b1),
    .dout(grp_fu_21385_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U43(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_18_fu_1441_p3),
    .din1(grp_fu_21397_p1),
    .ce(1'b1),
    .dout(grp_fu_21397_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U44(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21404_p0),
    .din1(grp_fu_21404_p1),
    .ce(1'b1),
    .dout(grp_fu_21404_p2)
);

mpc_mul_mul_21s_13s_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_13s_34_4_1_U45(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_19_fu_1589_p3),
    .din1(grp_fu_21411_p1),
    .ce(1'b1),
    .dout(grp_fu_21411_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U46(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21418_p0),
    .din1(grp_fu_21418_p1),
    .ce(1'b1),
    .dout(grp_fu_21418_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U47(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21430_p0),
    .din1(grp_fu_21430_p1),
    .ce(1'b1),
    .dout(grp_fu_21430_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U48(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21437_p0),
    .din1(grp_fu_21437_p1),
    .ce(1'b1),
    .dout(grp_fu_21437_p2)
);

mpc_mul_mul_21s_9s_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_9s_30_4_1_U49(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_5_fu_1741_p3),
    .din1(grp_fu_21449_p1),
    .ce(1'b1),
    .dout(grp_fu_21449_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U50(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_3_fu_1671_p3),
    .din1(grp_fu_21456_p1),
    .ce(1'b1),
    .dout(grp_fu_21456_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U51(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_5_fu_1741_p3),
    .din1(grp_fu_21465_p1),
    .ce(1'b1),
    .dout(grp_fu_21465_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U52(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_20_fu_1899_p3),
    .din1(grp_fu_21474_p1),
    .ce(1'b1),
    .dout(grp_fu_21474_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U53(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_7_fu_1969_p3),
    .din1(grp_fu_21481_p1),
    .ce(1'b1),
    .dout(grp_fu_21481_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U54(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21488_p0),
    .din1(grp_fu_21488_p1),
    .ce(1'b1),
    .dout(grp_fu_21488_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U55(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21495_p0),
    .din1(grp_fu_21495_p1),
    .ce(1'b1),
    .dout(grp_fu_21495_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U56(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_9_fu_2310_p3),
    .din1(grp_fu_21502_p1),
    .ce(1'b1),
    .dout(grp_fu_21502_p2)
);

mpc_mul_mul_21s_12ns_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_12ns_34_4_1_U57(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_10_fu_2993_p3),
    .din1(grp_fu_21509_p1),
    .ce(1'b1),
    .dout(grp_fu_21509_p2)
);

mpc_mul_mul_21s_8ns_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_8ns_30_4_1_U58(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_11_fu_3063_p3),
    .din1(grp_fu_21516_p1),
    .ce(1'b1),
    .dout(grp_fu_21516_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U59(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21523_p0),
    .din1(grp_fu_21523_p1),
    .ce(1'b1),
    .dout(grp_fu_21523_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U60(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21530_p0),
    .din1(grp_fu_21530_p1),
    .ce(1'b1),
    .dout(grp_fu_21530_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U61(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_11_fu_3063_p3),
    .din1(grp_fu_21539_p1),
    .ce(1'b1),
    .dout(grp_fu_21539_p2)
);

mpc_mul_mul_21s_15s_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_15s_36_4_1_U62(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_12_fu_3712_p3),
    .din1(grp_fu_21546_p1),
    .ce(1'b1),
    .dout(grp_fu_21546_p2)
);

mpc_mul_mul_21s_15s_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_15s_36_4_1_U63(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_13_fu_3782_p3),
    .din1(grp_fu_21553_p1),
    .ce(1'b1),
    .dout(grp_fu_21553_p2)
);

mpc_mul_mul_21s_14ns_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_14ns_36_4_1_U64(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_15_fu_4639_p3),
    .din1(grp_fu_21560_p1),
    .ce(1'b1),
    .dout(grp_fu_21560_p2)
);

mpc_mul_mul_21s_15s_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 15 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_15s_36_4_1_U65(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_14_fu_4569_p3),
    .din1(grp_fu_21567_p1),
    .ce(1'b1),
    .dout(grp_fu_21567_p2)
);

mpc_mul_mul_21s_14ns_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_14ns_36_4_1_U66(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_16_fu_5204_p3),
    .din1(grp_fu_21575_p1),
    .ce(1'b1),
    .dout(grp_fu_21575_p2)
);

mpc_mul_mul_21s_14ns_36_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 36 ))
mul_mul_21s_14ns_36_4_1_U67(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_17_fu_5274_p3),
    .din1(grp_fu_21582_p1),
    .ce(1'b1),
    .dout(grp_fu_21582_p2)
);

mpc_mul_mul_21s_9s_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_9s_30_4_1_U68(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21590_p0),
    .din1(grp_fu_21590_p1),
    .ce(1'b1),
    .dout(grp_fu_21590_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U69(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_23_fu_8709_p3),
    .din1(grp_fu_21597_p1),
    .ce(1'b1),
    .dout(grp_fu_21597_p2)
);

mpc_mul_mul_21s_10s_31_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 31 ))
mul_mul_21s_10s_31_4_1_U70(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_22_fu_9610_p3),
    .din1(grp_fu_21604_p1),
    .ce(1'b1),
    .dout(grp_fu_21604_p2)
);

mpc_mul_mul_21s_12ns_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_12ns_34_4_1_U71(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_22_fu_9610_p3),
    .din1(grp_fu_21611_p1),
    .ce(1'b1),
    .dout(grp_fu_21611_p2)
);

mpc_mul_mul_21s_12ns_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_12ns_34_4_1_U72(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_21_fu_10332_p3),
    .din1(grp_fu_21618_p1),
    .ce(1'b1),
    .dout(grp_fu_21618_p2)
);

mpc_mul_mul_21s_10s_31_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 10 ),
    .dout_WIDTH( 31 ))
mul_mul_21s_10s_31_4_1_U73(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_21_fu_10332_p3),
    .din1(grp_fu_21630_p1),
    .ce(1'b1),
    .dout(grp_fu_21630_p2)
);

mpc_mul_mul_21s_9s_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_9s_30_4_1_U74(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln302_21_fu_10332_p3),
    .din1(grp_fu_21642_p1),
    .ce(1'b1),
    .dout(grp_fu_21642_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U75(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21654_p0),
    .din1(grp_fu_21654_p1),
    .ce(1'b1),
    .dout(grp_fu_21654_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U76(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(select_ln346_139_fu_12187_p3),
    .din1(grp_fu_21666_p1),
    .ce(1'b1),
    .dout(grp_fu_21666_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U77(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21678_p0),
    .din1(grp_fu_21678_p1),
    .ce(1'b1),
    .dout(grp_fu_21678_p2)
);

mpc_mul_mul_21s_7ns_29_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 29 ))
mul_mul_21s_7ns_29_4_1_U78(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21690_p0),
    .din1(grp_fu_21690_p1),
    .ce(1'b1),
    .dout(grp_fu_21690_p2)
);

mpc_mul_mul_21s_12ns_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_12ns_34_4_1_U79(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21702_p0),
    .din1(grp_fu_21702_p1),
    .ce(1'b1),
    .dout(grp_fu_21702_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U80(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21714_p0),
    .din1(grp_fu_21714_p1),
    .ce(1'b1),
    .dout(grp_fu_21714_p2)
);

mpc_mul_mul_21s_8ns_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_8ns_30_4_1_U81(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21721_p0),
    .din1(grp_fu_21721_p1),
    .ce(1'b1),
    .dout(grp_fu_21721_p2)
);

mpc_mul_mul_21s_7ns_29_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 29 ))
mul_mul_21s_7ns_29_4_1_U82(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21733_p0),
    .din1(grp_fu_21733_p1),
    .ce(1'b1),
    .dout(grp_fu_21733_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U83(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21740_p0),
    .din1(grp_fu_21740_p1),
    .ce(1'b1),
    .dout(grp_fu_21740_p2)
);

mpc_mul_mul_21s_8s_29_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 29 ))
mul_mul_21s_8s_29_4_1_U84(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21752_p0),
    .din1(grp_fu_21752_p1),
    .ce(1'b1),
    .dout(grp_fu_21752_p2)
);

mpc_mul_mul_21s_13s_34_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 34 ))
mul_mul_21s_13s_34_4_1_U85(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21764_p0),
    .din1(grp_fu_21764_p1),
    .ce(1'b1),
    .dout(grp_fu_21764_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U86(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21776_p0),
    .din1(grp_fu_21776_p1),
    .ce(1'b1),
    .dout(grp_fu_21776_p2)
);

mpc_mul_mul_21s_9s_30_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 30 ))
mul_mul_21s_9s_30_4_1_U87(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21783_p0),
    .din1(grp_fu_21783_p1),
    .ce(1'b1),
    .dout(grp_fu_21783_p2)
);

mpc_mul_mul_21s_8s_29_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 8 ),
    .dout_WIDTH( 29 ))
mul_mul_21s_8s_29_4_1_U88(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21795_p0),
    .din1(grp_fu_21795_p1),
    .ce(1'b1),
    .dout(grp_fu_21795_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U89(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21802_p0),
    .din1(grp_fu_21802_p1),
    .ce(1'b1),
    .dout(grp_fu_21802_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U90(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21810_p0),
    .din1(grp_fu_21810_p1),
    .ce(1'b1),
    .dout(grp_fu_21810_p2)
);

mpc_mul_mul_21s_13ns_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_13ns_35_4_1_U91(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21819_p0),
    .din1(grp_fu_21819_p1),
    .ce(1'b1),
    .dout(grp_fu_21819_p2)
);

mpc_mul_mul_21s_6ns_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 6 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_6ns_28_4_1_U92(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21826_p0),
    .din1(grp_fu_21826_p1),
    .ce(1'b1),
    .dout(grp_fu_21826_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U93(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21833_p0),
    .din1(grp_fu_21833_p1),
    .ce(1'b1),
    .dout(grp_fu_21833_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U94(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21844_p0),
    .din1(grp_fu_21844_p1),
    .ce(1'b1),
    .dout(grp_fu_21844_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U95(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21855_p0),
    .din1(grp_fu_21855_p1),
    .ce(1'b1),
    .dout(grp_fu_21855_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U96(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21863_p0),
    .din1(grp_fu_21863_p1),
    .ce(1'b1),
    .dout(grp_fu_21863_p2)
);

mpc_mul_mul_21s_14s_35_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 14 ),
    .dout_WIDTH( 35 ))
mul_mul_21s_14s_35_4_1_U97(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21872_p0),
    .din1(grp_fu_21872_p1),
    .ce(1'b1),
    .dout(grp_fu_21872_p2)
);

mpc_mul_mul_21s_7s_28_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 21 ),
    .din1_WIDTH( 7 ),
    .dout_WIDTH( 28 ))
mul_mul_21s_7s_28_4_1_U98(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(grp_fu_21879_p0),
    .din1(grp_fu_21879_p1),
    .ce(1'b1),
    .dout(grp_fu_21879_p2)
);

mpc_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (ap_loop_exit_ready == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg <= 1'b0;
    end else begin
        if ((((1'b1 == ap_CS_fsm_state1) & (1'b1 == ap_NS_fsm_state2)) | ((1'b1 == ap_NS_fsm_state66) & (1'b1 == ap_CS_fsm_state65)) | ((1'b1 == ap_NS_fsm_state46) & (1'b1 == ap_CS_fsm_state45)) | ((1'b1 == ap_NS_fsm_state12) & (1'b1 == ap_CS_fsm_state11)))) begin
            grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg <= 1'b1;
        end else if ((grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_ready == 1'b1)) begin
            grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        if ((icmp_ln74_fu_1292_p2 == 1'd0)) begin
            i_fu_310 <= i_2_fu_1298_p2;
        end else if ((ap_loop_init == 1'b1)) begin
            i_fu_310 <= 5'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state27)) begin
        add_ln377_11_reg_23140 <= add_ln377_11_fu_9354_p2;
        and_ln895_46_reg_23145 <= and_ln895_46_fu_9456_p2;
        or_ln346_11_reg_23150 <= or_ln346_11_fu_9486_p2;
        select_ln302_22_reg_23155 <= select_ln302_22_fu_9610_p3;
        tmp_337_reg_23171 <= sub_ln1347_3_fu_9642_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state28)) begin
        add_ln377_12_reg_23176 <= add_ln377_12_fu_9715_p2;
        and_ln895_47_reg_23181 <= and_ln895_47_fu_9817_p2;
        mul_ln1273_28_reg_23191 <= grp_fu_21590_p2;
        mul_ln1273_32_reg_23202 <= grp_fu_21597_p2;
        or_ln346_12_reg_23186 <= or_ln346_12_fu_9847_p2;
        tmp_307_reg_23197 <= grp_fu_21590_p2[32'd13];
        tmp_343_reg_23208 <= grp_fu_21597_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state29)) begin
        add_ln377_13_reg_23213 <= add_ln377_13_fu_10026_p2;
        and_ln895_50_reg_23218 <= and_ln895_50_fu_10128_p2;
        or_ln346_13_reg_23223 <= or_ln346_13_fu_10158_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state18)) begin
        add_ln377_15_reg_22569 <= add_ln377_15_fu_3368_p2;
        add_ln377_25_reg_22605 <= add_ln377_25_fu_3542_p2;
        and_ln895_54_reg_22584 <= and_ln895_54_fu_3458_p2;
        and_ln895_70_reg_22620 <= and_ln895_70_fu_3632_p2;
        mul_ln1273_4_reg_22527 <= grp_fu_21449_p2;
        or_ln896_15_reg_22590 <= or_ln896_15_fu_3470_p2;
        or_ln896_25_reg_22626 <= or_ln896_25_fu_3644_p2;
        select_ln302_11_reg_22516 <= select_ln302_11_fu_3063_p3;
        select_ln346_40_reg_22522 <= select_ln346_40_fu_3271_p3;
        tmp_103_reg_22533 <= grp_fu_21449_p2[32'd13];
        tmp_169_reg_22559 <= add_ln1347_31_fu_3319_p2[32'd35];
        tmp_170_reg_22564 <= add_ln810_11_fu_3325_p2[32'd34];
        tmp_173_reg_22579 <= add_ln1347_31_fu_3319_p2[32'd35];
        tmp_241_reg_22595 <= add_ln1347_40_fu_3493_p2[32'd35];
        tmp_242_reg_22600 <= add_ln810_18_fu_3499_p2[32'd34];
        tmp_245_reg_22615 <= add_ln1347_40_fu_3493_p2[32'd35];
        xor_ln896_34_reg_22574 <= xor_ln896_34_fu_3382_p2;
        xor_ln896_60_reg_22610 <= xor_ln896_60_fu_3556_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state19)) begin
        add_ln377_16_reg_22673 <= add_ln377_16_fu_4127_p2;
        add_ln377_3_reg_22631 <= add_ln377_3_fu_3878_p2;
        and_ln895_38_reg_22636 <= and_ln895_38_fu_3980_p2;
        and_ln895_55_reg_22678 <= and_ln895_55_fu_4229_p2;
        mul_ln1273_5_reg_22646 <= grp_fu_21474_p2;
        mul_ln1273_6_reg_22657 <= grp_fu_21481_p2;
        or_ln346_16_reg_22683 <= or_ln346_16_fu_4259_p2;
        or_ln346_3_reg_22641 <= or_ln346_3_fu_4010_p2;
        select_ln346_114_reg_22693 <= select_ln346_114_fu_4499_p3;
        tmp_109_reg_22652 <= grp_fu_21474_p2[32'd13];
        tmp_115_reg_22663 <= grp_fu_21481_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state20)) begin
        add_ln377_17_reg_22719 <= add_ln377_17_fu_4986_p2;
        and_ln895_56_reg_22724 <= and_ln895_56_fu_5088_p2;
        mul_ln1273_15_reg_22734 <= grp_fu_21495_p2;
        mul_ln1273_16_reg_22745 <= grp_fu_21502_p2;
        mul_ln1273_7_reg_22703 <= grp_fu_21488_p2;
        or_ln346_17_reg_22729 <= or_ln346_17_fu_5118_p2;
        select_ln346_44_reg_22698 <= select_ln346_44_fu_4865_p3;
        tmp_121_reg_22709 <= grp_fu_21488_p2[32'd13];
        tmp_193_reg_22740 <= grp_fu_21495_p2[32'd13];
        tmp_199_reg_22751 <= grp_fu_21502_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state21)) begin
        add_ln377_18_reg_22798 <= add_ln377_18_fu_5676_p2;
        add_ln377_26_reg_22850 <= add_ln377_26_fu_5857_p2;
        and_ln895_59_reg_22813 <= and_ln895_59_fu_5766_p2;
        and_ln895_75_reg_22865 <= and_ln895_75_fu_5947_p2;
        mul_ln1273_17_reg_22824 <= grp_fu_21523_p2;
        mul_ln1273_23_reg_22876 <= grp_fu_21539_p2;
        mul_ln1273_8_reg_22766 <= grp_fu_21509_p2;
        mul_ln1273_9_reg_22777 <= grp_fu_21516_p2;
        or_ln896_18_reg_22819 <= or_ln896_18_fu_5778_p2;
        or_ln896_26_reg_22871 <= or_ln896_26_fu_5959_p2;
        select_ln346_46_reg_22761 <= select_ln346_46_fu_5486_p3;
        tmp_133_reg_22772 <= grp_fu_21509_p2[32'd13];
        tmp_139_reg_22783 <= grp_fu_21516_p2[32'd13];
        tmp_191_reg_22788 <= add_ln1347_34_fu_5636_p2[32'd35];
        tmp_192_reg_22793 <= add_ln810_14_fu_5642_p2[32'd34];
        tmp_195_reg_22808 <= add_ln1347_34_fu_5636_p2[32'd35];
        tmp_205_reg_22830 <= grp_fu_21523_p2[32'd13];
        tmp_255_reg_22840 <= add_ln1347_41_fu_5809_p2[32'd35];
        tmp_256_reg_22845 <= add_ln810_19_fu_5815_p2[32'd34];
        tmp_259_reg_22860 <= add_ln1347_41_fu_5809_p2[32'd35];
        tmp_263_reg_22882 <= grp_fu_21539_p2[32'd13];
        xor_ln896_42_reg_22803 <= xor_ln896_42_fu_5690_p2;
        xor_ln896_66_reg_22855 <= xor_ln896_66_fu_5871_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state22)) begin
        add_ln377_19_reg_22907 <= add_ln377_19_fu_6288_p2;
        add_ln377_27_reg_22932 <= add_ln377_27_fu_6530_p2;
        and_ln895_60_reg_22912 <= and_ln895_60_fu_6390_p2;
        and_ln895_76_reg_22937 <= and_ln895_76_fu_6632_p2;
        mul_ln1273_10_reg_22897 <= grp_fu_21546_p2;
        mul_ln1273_18_reg_22922 <= grp_fu_21553_p2;
        or_ln346_19_reg_22917 <= or_ln346_19_fu_6420_p2;
        or_ln346_27_reg_22942 <= or_ln346_27_fu_6662_p2;
        select_ln346_48_reg_22892 <= select_ln346_48_fu_6176_p3;
        tmp_145_reg_22902 <= grp_fu_21546_p2[32'd13];
        tmp_219_reg_22927 <= grp_fu_21553_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state24)) begin
        add_ln377_21_reg_23008 <= add_ln377_21_fu_7689_p2;
        add_ln377_29_reg_23043 <= add_ln377_29_fu_8026_p2;
        and_ln895_62_reg_23013 <= and_ln895_62_fu_7791_p2;
        and_ln895_82_reg_23058 <= and_ln895_82_fu_8116_p2;
        mul_ln1273_19_reg_23023 <= grp_fu_21575_p2;
        or_ln346_21_reg_23018 <= or_ln346_21_fu_7821_p2;
        or_ln896_29_reg_23064 <= or_ln896_29_fu_8128_p2;
        select_ln346_52_reg_23003 <= select_ln346_52_fu_7584_p3;
        tmp_229_reg_23028 <= grp_fu_21575_p2[32'd13];
        tmp_281_reg_23033 <= add_ln1347_44_fu_7984_p2[32'd35];
        tmp_282_reg_23038 <= add_ln1347_44_fu_7984_p2[32'd34];
        tmp_285_reg_23053 <= add_ln1347_44_fu_7984_p2[32'd35];
        xor_ln896_76_reg_23048 <= xor_ln896_76_fu_8040_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        add_ln377_22_reg_23084 <= add_ln377_22_fu_8478_p2;
        add_ln377_9_reg_23069 <= add_ln377_9_fu_8231_p2;
        and_ln895_44_reg_23074 <= and_ln895_44_fu_8333_p2;
        and_ln895_64_reg_23089 <= and_ln895_64_fu_8580_p2;
        or_ln346_22_reg_23094 <= or_ln346_22_fu_8610_p2;
        or_ln346_9_reg_23079 <= or_ln346_9_fu_8363_p2;
        sub_ln1273_4_reg_23109 <= sub_ln1273_4_fu_8753_p2;
        tmp_325_reg_23115 <= sub_ln1347_2_fu_8759_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state26)) begin
        add_ln377_23_reg_23125 <= add_ln377_23_fu_9158_p2;
        and_ln895_67_reg_23130 <= and_ln895_67_fu_9260_p2;
        or_ln346_23_reg_23135 <= or_ln346_23_fu_9290_p2;
        select_ln346_56_reg_23120 <= select_ln346_56_fu_8991_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state23)) begin
        add_ln377_28_reg_22977 <= add_ln377_28_fu_7276_p2;
        and_ln895_79_reg_22992 <= and_ln895_79_fu_7366_p2;
        mul_ln1273_11_reg_22952 <= grp_fu_21560_p2;
        or_ln896_28_reg_22998 <= or_ln896_28_fu_7378_p2;
        select_ln346_50_reg_22947 <= select_ln346_50_fu_6872_p3;
        select_ln346_88_reg_22962 <= select_ln346_88_fu_7101_p3;
        tmp_155_reg_22957 <= grp_fu_21560_p2[32'd13];
        tmp_271_reg_22967 <= add_ln1347_43_fu_7234_p2[32'd35];
        tmp_272_reg_22972 <= add_ln1347_43_fu_7234_p2[32'd34];
        tmp_275_reg_22987 <= add_ln1347_43_fu_7234_p2[32'd35];
        xor_ln896_72_reg_22982 <= xor_ln896_72_fu_7290_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state35)) begin
        add_ln377_32_reg_23325 <= add_ln377_32_fu_11640_p2;
        add_ln377_35_reg_23340 <= add_ln377_35_fu_11836_p2;
        add_ln377_38_reg_23355 <= add_ln377_38_fu_12042_p2;
        and_ln895_88_reg_23330 <= and_ln895_88_fu_11742_p2;
        and_ln895_91_reg_23345 <= and_ln895_91_fu_11938_p2;
        and_ln895_94_reg_23360 <= and_ln895_94_fu_12144_p2;
        or_ln346_32_reg_23335 <= or_ln346_32_fu_11772_p2;
        or_ln346_35_reg_23350 <= or_ln346_35_fu_11968_p2;
        or_ln346_38_reg_23365 <= or_ln346_38_fu_12174_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state33)) begin
        add_ln377_33_reg_23270 <= add_ln377_33_fu_10594_p2;
        add_ln377_36_reg_23285 <= add_ln377_36_fu_10768_p2;
        and_ln895_89_reg_23275 <= and_ln895_89_fu_10694_p2;
        and_ln895_92_reg_23290 <= and_ln895_92_fu_10868_p2;
        or_ln346_33_reg_23280 <= or_ln346_33_fu_10724_p2;
        or_ln346_36_reg_23295 <= or_ln346_36_fu_10898_p2;
        select_ln346_135_reg_23265 <= select_ln346_135_fu_10548_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state34)) begin
        add_ln377_37_reg_23310 <= add_ln377_37_fu_11444_p2;
        and_ln895_93_reg_23315 <= and_ln895_93_fu_11546_p2;
        or_ln346_37_reg_23320 <= or_ln346_37_fu_11576_p2;
        select_ln346_137_reg_23300 <= select_ln346_137_fu_11111_p3;
        select_ln346_143_reg_23305 <= select_ln346_143_fu_11341_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state39)) begin
        add_ln377_39_reg_23450 <= add_ln377_39_fu_13145_p2;
        add_ln377_40_reg_23465 <= add_ln377_40_fu_13319_p2;
        add_ln377_43_reg_23485 <= add_ln377_43_fu_13679_p2;
        add_ln377_48_reg_23516 <= add_ln377_48_fu_14050_p2;
        add_ln377_55_reg_23547 <= add_ln377_55_fu_14417_p2;
        add_ln377_60_reg_23578 <= add_ln377_60_fu_14788_p2;
        and_ln895_104_reg_23490 <= and_ln895_104_fu_13779_p2;
        and_ln895_110_reg_23521 <= and_ln895_110_fu_14150_p2;
        and_ln895_122_reg_23552 <= and_ln895_122_fu_14517_p2;
        and_ln895_128_reg_23583 <= and_ln895_128_fu_14888_p2;
        and_ln895_95_reg_23455 <= and_ln895_95_fu_13245_p2;
        and_ln895_98_reg_23470 <= and_ln895_98_fu_13419_p2;
        mul_ln1273_40_reg_23500 <= grp_fu_21714_p2;
        mul_ln1273_43_reg_23531 <= grp_fu_21733_p2;
        mul_ln1273_52_reg_23562 <= grp_fu_21776_p2;
        mul_ln1273_55_reg_23593 <= grp_fu_21795_p2;
        or_ln346_39_reg_23460 <= or_ln346_39_fu_13275_p2;
        or_ln346_40_reg_23475 <= or_ln346_40_fu_13449_p2;
        or_ln346_43_reg_23495 <= or_ln346_43_fu_13809_p2;
        or_ln346_48_reg_23526 <= or_ln346_48_fu_14180_p2;
        or_ln346_55_reg_23557 <= or_ln346_55_fu_14547_p2;
        or_ln346_60_reg_23588 <= or_ln346_60_fu_14918_p2;
        select_ln346_165_reg_23480 <= select_ln346_165_fu_13633_p3;
        select_ln346_177_reg_23506 <= select_ln346_177_fu_13997_p3;
        select_ln346_201_reg_23542 <= select_ln346_201_fu_14371_p3;
        select_ln346_213_reg_23568 <= select_ln346_213_fu_14735_p3;
        tmp_403_reg_23511 <= grp_fu_21714_p2[32'd13];
        tmp_421_reg_23537 <= grp_fu_21733_p2[32'd13];
        tmp_487_reg_23573 <= grp_fu_21776_p2[32'd13];
        tmp_505_reg_23599 <= grp_fu_21795_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state40)) begin
        add_ln377_42_reg_23614 <= add_ln377_42_fu_15225_p2;
        add_ln377_44_reg_23650 <= add_ln377_44_fu_15417_p2;
        add_ln377_51_reg_23708 <= add_ln377_51_fu_16011_p2;
        add_ln377_52_reg_23723 <= add_ln377_52_fu_16185_p2;
        add_ln377_54_reg_23748 <= add_ln377_54_fu_16383_p2;
        add_ln377_56_reg_23784 <= add_ln377_56_fu_16575_p2;
        and_ln895_102_reg_23629 <= and_ln895_102_fu_15315_p2;
        and_ln895_105_reg_23665 <= and_ln895_105_fu_15507_p2;
        and_ln895_113_reg_23713 <= and_ln895_113_fu_16111_p2;
        and_ln895_116_reg_23728 <= and_ln895_116_fu_16285_p2;
        and_ln895_120_reg_23763 <= and_ln895_120_fu_16473_p2;
        and_ln895_123_reg_23799 <= and_ln895_123_fu_16665_p2;
        mul_ln1273_41_reg_23676 <= grp_fu_21819_p2;
        mul_ln1273_44_reg_23692 <= grp_fu_21826_p2;
        mul_ln1273_53_reg_23810 <= grp_fu_21872_p2;
        mul_ln1273_56_reg_23826 <= grp_fu_21879_p2;
        or_ln346_51_reg_23718 <= or_ln346_51_fu_16141_p2;
        or_ln346_52_reg_23733 <= or_ln346_52_fu_16315_p2;
        or_ln896_42_reg_23635 <= or_ln896_42_fu_15327_p2;
        or_ln896_44_reg_23671 <= or_ln896_44_fu_15519_p2;
        or_ln896_54_reg_23769 <= or_ln896_54_fu_16485_p2;
        or_ln896_56_reg_23805 <= or_ln896_56_fu_16677_p2;
        select_ln346_179_reg_23682 <= select_ln346_179_fu_15725_p3;
        select_ln346_185_reg_23698 <= select_ln346_185_fu_15962_p3;
        select_ln346_215_reg_23816 <= select_ln346_215_fu_16883_p3;
        select_ln346_221_reg_23832 <= select_ln346_221_fu_17120_p3;
        tmp_373_reg_23604 <= add_ln1347_51_fu_15177_p2[32'd35];
        tmp_374_reg_23609 <= add_ln810_27_fu_15183_p2[32'd34];
        tmp_377_reg_23624 <= add_ln1347_51_fu_15177_p2[32'd35];
        tmp_387_reg_23640 <= add_ln1347_52_fu_15368_p2[32'd35];
        tmp_388_reg_23645 <= add_ln810_28_fu_15374_p2[32'd34];
        tmp_391_reg_23660 <= add_ln1347_52_fu_15368_p2[32'd35];
        tmp_409_reg_23687 <= grp_fu_21819_p2[32'd13];
        tmp_427_reg_23703 <= grp_fu_21826_p2[32'd13];
        tmp_457_reg_23738 <= add_ln1347_57_fu_16335_p2[32'd35];
        tmp_458_reg_23743 <= add_ln810_33_fu_16341_p2[32'd34];
        tmp_461_reg_23758 <= add_ln1347_57_fu_16335_p2[32'd35];
        tmp_471_reg_23774 <= add_ln1347_58_fu_16526_p2[32'd35];
        tmp_472_reg_23779 <= add_ln810_34_fu_16532_p2[32'd34];
        tmp_475_reg_23794 <= add_ln1347_58_fu_16526_p2[32'd35];
        tmp_493_reg_23821 <= grp_fu_21872_p2[32'd13];
        tmp_511_reg_23837 <= grp_fu_21879_p2[32'd13];
        xor_ln896_106_reg_23619 <= xor_ln896_106_fu_15239_p2;
        xor_ln896_111_reg_23655 <= xor_ln896_111_fu_15431_p2;
        xor_ln896_136_reg_23753 <= xor_ln896_136_fu_16397_p2;
        xor_ln896_141_reg_23789 <= xor_ln896_141_fu_16589_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        mul_ln1273_14_reg_22500 <= grp_fu_21430_p2;
        mul_ln1273_2_reg_22457 <= grp_fu_21404_p2;
        mul_ln1273_3_reg_22473 <= grp_fu_21411_p2;
        select_ln302_9_reg_22451 <= select_ln302_9_fu_2310_p3;
        select_ln346_104_reg_22511 <= select_ln346_104_fu_2923_p3;
        select_ln346_38_reg_22463 <= select_ln346_38_fu_2522_p3;
        select_ln346_72_reg_22495 <= select_ln346_72_fu_2730_p3;
        tmp_177_reg_22506 <= grp_fu_21430_p2[32'd13];
        tmp_85_reg_22468 <= grp_fu_21404_p2[32'd13];
        tmp_97_reg_22479 <= grp_fu_21411_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state16)) begin
        mul_ln1273_1_reg_22425 <= grp_fu_21397_p2;
        select_ln346_36_reg_22431 <= select_ln346_36_fu_2155_p3;
        tmp_79_reg_22436 <= grp_fu_21397_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state30)) begin
        mul_ln1273_27_reg_23243 <= grp_fu_21604_p2;
        mul_ln1273_30_reg_23254 <= grp_fu_21611_p2;
        tmp_301_reg_23249 <= grp_fu_21604_p2[32'd13];
        tmp_319_reg_23260 <= grp_fu_21611_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state2))) begin
        reg_1200 <= uk_admm_V_q1;
        reg_1204 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state3))) begin
        reg_1208 <= uk_admm_V_q1;
        reg_1212 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state4))) begin
        reg_1216 <= uk_admm_V_q1;
        reg_1220 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state5))) begin
        reg_1224 <= uk_admm_V_q1;
        reg_1228 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state6))) begin
        reg_1232 <= uk_admm_V_q1;
        reg_1236 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state7))) begin
        reg_1240 <= uk_admm_V_q1;
        reg_1244 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state8))) begin
        reg_1248 <= uk_admm_V_q1;
        reg_1252 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state9))) begin
        reg_1256 <= uk_admm_V_q1;
        reg_1260 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state10))) begin
        reg_1264 <= uk_admm_V_q1;
        reg_1268 <= uk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state15)) begin
        select_ln302_3_reg_22388 <= select_ln302_3_fu_1671_p3;
        select_ln302_5_reg_22394 <= select_ln302_5_fu_1741_p3;
        tmp_183_reg_22420 <= sub_ln1347_1_fu_1823_p2[32'd13];
        tmp_91_reg_22405 <= sub_ln1347_fu_1777_p2[32'd13];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state36)) begin
        select_ln346_139_reg_23370 <= select_ln346_139_fu_12187_p3;
        select_ln346_145_reg_23375 <= select_ln346_145_fu_12206_p3;
        sext_ln1273_43_reg_23399 <= sext_ln1273_43_fu_12224_p1;
        sext_ln1273_44_reg_23405 <= sext_ln1273_44_fu_12228_p1;
        sext_ln1273_47_reg_23419 <= sext_ln1273_47_fu_12236_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state37)) begin
        select_ln346_151_reg_23427 <= select_ln346_151_fu_12531_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state41)) begin
        select_ln346_169_reg_23842 <= select_ln346_169_fu_17215_p3;
        select_ln346_175_reg_23847 <= select_ln346_175_fu_17303_p3;
        select_ln346_181_reg_23852 <= select_ln346_181_fu_17511_p3;
        select_ln346_187_reg_23857 <= select_ln346_187_fu_17723_p3;
        select_ln346_205_reg_23862 <= select_ln346_205_fu_18043_p3;
        select_ln346_211_reg_23867 <= select_ln346_211_fu_18131_p3;
        select_ln346_217_reg_23872 <= select_ln346_217_fu_18339_p3;
        select_ln346_223_reg_23877 <= select_ln346_223_fu_18551_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        sext_ln813_71_reg_21983 <= sext_ln813_71_fu_1272_p1;
        sext_ln813_72_reg_21988 <= sext_ln813_72_fu_1276_p1;
        sext_ln813_73_reg_21993 <= sext_ln813_73_fu_1280_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state72)) begin
        zk_admm_V_load_10_reg_23942 <= zk_admm_V_q1;
        zk_admm_V_load_11_reg_23948 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state73)) begin
        zk_admm_V_load_12_reg_23954 <= zk_admm_V_q1;
        zk_admm_V_load_13_reg_23960 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state74)) begin
        zk_admm_V_load_14_reg_23966 <= zk_admm_V_q1;
        zk_admm_V_load_15_reg_23972 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state75)) begin
        zk_admm_V_load_16_reg_23978 <= zk_admm_V_q1;
        zk_admm_V_load_17_reg_23984 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state67)) begin
        zk_admm_V_load_1_reg_23888 <= zk_admm_V_q0;
        zk_admm_V_load_reg_23882 <= zk_admm_V_q1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state68)) begin
        zk_admm_V_load_2_reg_23894 <= zk_admm_V_q1;
        zk_admm_V_load_3_reg_23900 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state69)) begin
        zk_admm_V_load_4_reg_23906 <= zk_admm_V_q1;
        zk_admm_V_load_5_reg_23912 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state70)) begin
        zk_admm_V_load_6_reg_23918 <= zk_admm_V_q1;
        zk_admm_V_load_7_reg_23924 <= zk_admm_V_q0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state71)) begin
        zk_admm_V_load_8_reg_23930 <= zk_admm_V_q1;
        zk_admm_V_load_9_reg_23936 <= zk_admm_V_q0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state45))) begin
        Hxk_V_address0 = 64'd11;
    end else if (((1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state44))) begin
        Hxk_V_address0 = 64'd5;
    end else if (((1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state43))) begin
        Hxk_V_address0 = 64'd9;
    end else if (((1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state42))) begin
        Hxk_V_address0 = 64'd3;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state41))) begin
        Hxk_V_address0 = 64'd7;
    end else if (((1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_address0 = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state38))) begin
        Hxk_V_address0 = 64'd17;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state63))) begin
        Hxk_V_address0 = 64'd15;
    end else if (((1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state62))) begin
        Hxk_V_address0 = 64'd13;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        Hxk_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address0;
    end else begin
        Hxk_V_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state45))) begin
        Hxk_V_address1 = 64'd10;
    end else if (((1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state44))) begin
        Hxk_V_address1 = 64'd4;
    end else if (((1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state43))) begin
        Hxk_V_address1 = 64'd8;
    end else if (((1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state42))) begin
        Hxk_V_address1 = 64'd2;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state41))) begin
        Hxk_V_address1 = 64'd6;
    end else if (((1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_address1 = 64'd0;
    end else if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state38))) begin
        Hxk_V_address1 = 64'd16;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state63))) begin
        Hxk_V_address1 = 64'd14;
    end else if (((1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state62))) begin
        Hxk_V_address1 = 64'd12;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        Hxk_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address1;
    end else begin
        Hxk_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state45) | (1'b1 == ap_CS_fsm_state41) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        Hxk_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce0;
    end else begin
        Hxk_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state45) | (1'b1 == ap_CS_fsm_state41) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        Hxk_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce1;
    end else begin
        Hxk_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state45)) begin
        Hxk_V_d0 = select_ln346_223_reg_23877;
    end else if ((1'b1 == ap_CS_fsm_state44)) begin
        Hxk_V_d0 = select_ln346_187_reg_23857;
    end else if ((1'b1 == ap_CS_fsm_state43)) begin
        Hxk_V_d0 = select_ln346_211_reg_23867;
    end else if ((1'b1 == ap_CS_fsm_state42)) begin
        Hxk_V_d0 = select_ln346_175_reg_23847;
    end else if ((1'b1 == ap_CS_fsm_state41)) begin
        Hxk_V_d0 = select_ln346_199_fu_17954_p3;
    end else if ((1'b1 == ap_CS_fsm_state40)) begin
        Hxk_V_d0 = select_ln346_163_fu_15154_p3;
    end else if ((1'b1 == ap_CS_fsm_state38)) begin
        Hxk_V_d0 = select_ln346_247_fu_13102_p3;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        Hxk_V_d0 = select_ln346_241_fu_12832_p3;
    end else if ((1'b1 == ap_CS_fsm_state36)) begin
        Hxk_V_d0 = select_ln346_233_fu_12515_p3;
    end else begin
        Hxk_V_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state45)) begin
        Hxk_V_d1 = select_ln346_217_reg_23872;
    end else if ((1'b1 == ap_CS_fsm_state44)) begin
        Hxk_V_d1 = select_ln346_181_reg_23852;
    end else if ((1'b1 == ap_CS_fsm_state43)) begin
        Hxk_V_d1 = select_ln346_205_reg_23862;
    end else if ((1'b1 == ap_CS_fsm_state42)) begin
        Hxk_V_d1 = select_ln346_169_reg_23842;
    end else if ((1'b1 == ap_CS_fsm_state41)) begin
        Hxk_V_d1 = select_ln346_193_fu_17836_p3;
    end else if ((1'b1 == ap_CS_fsm_state40)) begin
        Hxk_V_d1 = select_ln346_157_fu_15036_p3;
    end else if ((1'b1 == ap_CS_fsm_state38)) begin
        Hxk_V_d1 = select_ln346_245_fu_13003_p3;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        Hxk_V_d1 = select_ln346_235_fu_12622_p3;
    end else if ((1'b1 == ap_CS_fsm_state36)) begin
        Hxk_V_d1 = select_ln346_229_fu_12382_p3;
    end else begin
        Hxk_V_d1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state45) | (1'b1 == ap_CS_fsm_state41) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_we0 = 1'b1;
    end else begin
        Hxk_V_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state45) | (1'b1 == ap_CS_fsm_state41) | (1'b1 == ap_CS_fsm_state40))) begin
        Hxk_V_we1 = 1'b1;
    end else begin
        Hxk_V_we1 = 1'b0;
    end
end

assign ap_ST_fsm_state10_blk = 1'b0;

assign ap_ST_fsm_state11_blk = 1'b0;

assign ap_ST_fsm_state12_blk = 1'b0;

assign ap_ST_fsm_state13_blk = 1'b0;

assign ap_ST_fsm_state14_blk = 1'b0;

assign ap_ST_fsm_state15_blk = 1'b0;

assign ap_ST_fsm_state16_blk = 1'b0;

assign ap_ST_fsm_state17_blk = 1'b0;

assign ap_ST_fsm_state18_blk = 1'b0;

assign ap_ST_fsm_state19_blk = 1'b0;

always @ (*) begin
    if ((ap_start_int == 1'b0)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

assign ap_ST_fsm_state20_blk = 1'b0;

assign ap_ST_fsm_state21_blk = 1'b0;

assign ap_ST_fsm_state22_blk = 1'b0;

assign ap_ST_fsm_state23_blk = 1'b0;

assign ap_ST_fsm_state24_blk = 1'b0;

assign ap_ST_fsm_state25_blk = 1'b0;

assign ap_ST_fsm_state26_blk = 1'b0;

assign ap_ST_fsm_state27_blk = 1'b0;

assign ap_ST_fsm_state28_blk = 1'b0;

assign ap_ST_fsm_state29_blk = 1'b0;

assign ap_ST_fsm_state2_blk = 1'b0;

assign ap_ST_fsm_state30_blk = 1'b0;

assign ap_ST_fsm_state31_blk = 1'b0;

assign ap_ST_fsm_state32_blk = 1'b0;

assign ap_ST_fsm_state33_blk = 1'b0;

assign ap_ST_fsm_state34_blk = 1'b0;

assign ap_ST_fsm_state35_blk = 1'b0;

assign ap_ST_fsm_state36_blk = 1'b0;

assign ap_ST_fsm_state37_blk = 1'b0;

assign ap_ST_fsm_state38_blk = 1'b0;

assign ap_ST_fsm_state39_blk = 1'b0;

assign ap_ST_fsm_state3_blk = 1'b0;

assign ap_ST_fsm_state40_blk = 1'b0;

assign ap_ST_fsm_state41_blk = 1'b0;

assign ap_ST_fsm_state42_blk = 1'b0;

assign ap_ST_fsm_state43_blk = 1'b0;

assign ap_ST_fsm_state44_blk = 1'b0;

assign ap_ST_fsm_state45_blk = 1'b0;

assign ap_ST_fsm_state46_blk = 1'b0;

assign ap_ST_fsm_state47_blk = 1'b0;

assign ap_ST_fsm_state48_blk = 1'b0;

assign ap_ST_fsm_state49_blk = 1'b0;

assign ap_ST_fsm_state4_blk = 1'b0;

assign ap_ST_fsm_state50_blk = 1'b0;

assign ap_ST_fsm_state51_blk = 1'b0;

assign ap_ST_fsm_state52_blk = 1'b0;

assign ap_ST_fsm_state53_blk = 1'b0;

assign ap_ST_fsm_state54_blk = 1'b0;

assign ap_ST_fsm_state55_blk = 1'b0;

assign ap_ST_fsm_state56_blk = 1'b0;

assign ap_ST_fsm_state57_blk = 1'b0;

assign ap_ST_fsm_state58_blk = 1'b0;

assign ap_ST_fsm_state59_blk = 1'b0;

assign ap_ST_fsm_state5_blk = 1'b0;

assign ap_ST_fsm_state60_blk = 1'b0;

assign ap_ST_fsm_state61_blk = 1'b0;

assign ap_ST_fsm_state62_blk = 1'b0;

assign ap_ST_fsm_state63_blk = 1'b0;

assign ap_ST_fsm_state64_blk = 1'b0;

assign ap_ST_fsm_state65_blk = 1'b0;

assign ap_ST_fsm_state66_blk = 1'b0;

assign ap_ST_fsm_state67_blk = 1'b0;

assign ap_ST_fsm_state68_blk = 1'b0;

assign ap_ST_fsm_state69_blk = 1'b0;

assign ap_ST_fsm_state6_blk = 1'b0;

assign ap_ST_fsm_state70_blk = 1'b0;

assign ap_ST_fsm_state71_blk = 1'b0;

assign ap_ST_fsm_state72_blk = 1'b0;

assign ap_ST_fsm_state73_blk = 1'b0;

assign ap_ST_fsm_state74_blk = 1'b0;

assign ap_ST_fsm_state75_blk = 1'b0;

assign ap_ST_fsm_state76_blk = 1'b0;

assign ap_ST_fsm_state77_blk = 1'b0;

assign ap_ST_fsm_state78_blk = 1'b0;

assign ap_ST_fsm_state79_blk = 1'b0;

assign ap_ST_fsm_state7_blk = 1'b0;

assign ap_ST_fsm_state80_blk = 1'b0;

assign ap_ST_fsm_state81_blk = 1'b0;

assign ap_ST_fsm_state82_blk = 1'b0;

assign ap_ST_fsm_state83_blk = 1'b0;

assign ap_ST_fsm_state84_blk = 1'b0;

assign ap_ST_fsm_state85_blk = 1'b0;

assign ap_ST_fsm_state8_blk = 1'b0;

assign ap_ST_fsm_state9_blk = 1'b0;

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (icmp_ln74_fu_1292_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter0_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter0_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (ap_loop_exit_ready == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state85)) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_loop_init == 1'b1))) begin
        ap_sig_allocacmp_i_1 = 5'd0;
    end else begin
        ap_sig_allocacmp_i_1 = i_fu_310;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0 = temp6_V_q0;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0 = temp4_V_q0;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0 = h_q0;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0 = zk_admm_V_q0;
    end else begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1 = temp6_V_q1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1 = temp4_V_q1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1 = h_q1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1 = zk_admm_V_q1;
    end else begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_q1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0 = Hxk_V_q0;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0 = uk_admm_V_q0;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0 = h_q0;
    end else begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1 = Hxk_V_q1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1 = uk_admm_V_q1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1 = h_q1;
    end else begin
        grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_q1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        h_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address0;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        h_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0;
    end else begin
        h_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        h_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        h_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1;
    end else begin
        h_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        h_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce0;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        h_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0;
    end else begin
        h_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        h_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        h_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1;
    end else begin
        h_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        temp4_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0;
    end else begin
        temp4_V_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        temp4_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1;
    end else begin
        temp4_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        temp4_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0;
    end else begin
        temp4_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state46))) begin
        temp4_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1;
    end else begin
        temp4_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_we0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0;
    end else begin
        temp4_V_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13))) begin
        temp4_V_we1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1;
    end else begin
        temp4_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state64)) begin
        temp5_address0 = 64'd17;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp5_address0 = 64'd15;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp5_address0 = 64'd13;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp5_address0 = 64'd11;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp5_address0 = 64'd9;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp5_address0 = 64'd7;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp5_address0 = 64'd5;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp5_address0 = 64'd3;
    end else if ((1'b1 == ap_CS_fsm_state56)) begin
        temp5_address0 = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0;
    end else begin
        temp5_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state64)) begin
        temp5_address1 = 64'd16;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp5_address1 = 64'd14;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp5_address1 = 64'd12;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp5_address1 = 64'd10;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp5_address1 = 64'd8;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp5_address1 = 64'd6;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp5_address1 = 64'd4;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp5_address1 = 64'd2;
    end else if ((1'b1 == ap_CS_fsm_state56)) begin
        temp5_address1 = 64'd0;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1;
    end else begin
        temp5_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state56))) begin
        temp5_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0;
    end else begin
        temp5_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state56))) begin
        temp5_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1;
    end else begin
        temp5_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_we0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0;
    end else begin
        temp5_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state49) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state47))) begin
        temp5_we1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1;
    end else begin
        temp5_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        temp6_V_address0 = 64'd17;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        temp6_V_address0 = 64'd15;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp6_V_address0 = 64'd13;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp6_V_address0 = 64'd11;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp6_V_address0 = 64'd9;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp6_V_address0 = 64'd7;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp6_V_address0 = 64'd5;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp6_V_address0 = 64'd3;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp6_V_address0 = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp6_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0;
    end else begin
        temp6_V_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        temp6_V_address1 = 64'd16;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        temp6_V_address1 = 64'd14;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp6_V_address1 = 64'd12;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp6_V_address1 = 64'd10;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp6_V_address1 = 64'd8;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp6_V_address1 = 64'd6;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp6_V_address1 = 64'd4;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp6_V_address1 = 64'd2;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp6_V_address1 = 64'd0;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp6_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1;
    end else begin
        temp6_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        temp6_V_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp6_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0;
    end else begin
        temp6_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        temp6_V_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp6_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1;
    end else begin
        temp6_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        temp6_V_d0 = select_ln302_41_fu_20100_p3;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        temp6_V_d0 = select_ln302_39_fu_19924_p3;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp6_V_d0 = select_ln302_37_fu_19748_p3;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp6_V_d0 = select_ln302_35_fu_19572_p3;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp6_V_d0 = select_ln302_33_fu_19396_p3;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp6_V_d0 = select_ln302_31_fu_19220_p3;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp6_V_d0 = select_ln302_29_fu_19044_p3;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp6_V_d0 = select_ln302_27_fu_18868_p3;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp6_V_d0 = select_ln302_25_fu_18692_p3;
    end else begin
        temp6_V_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        temp6_V_d1 = select_ln302_40_fu_20029_p3;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        temp6_V_d1 = select_ln302_38_fu_19853_p3;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        temp6_V_d1 = select_ln302_36_fu_19677_p3;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        temp6_V_d1 = select_ln302_34_fu_19501_p3;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        temp6_V_d1 = select_ln302_32_fu_19325_p3;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        temp6_V_d1 = select_ln302_30_fu_19149_p3;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        temp6_V_d1 = select_ln302_28_fu_18973_p3;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        temp6_V_d1 = select_ln302_26_fu_18797_p3;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        temp6_V_d1 = select_ln302_24_fu_18621_p3;
    end else begin
        temp6_V_d1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        temp6_V_we0 = 1'b1;
    end else begin
        temp6_V_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        temp6_V_we1 = 1'b1;
    end else begin
        temp6_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state84)) begin
        temp7_address0 = 64'd17;
    end else if ((1'b1 == ap_CS_fsm_state83)) begin
        temp7_address0 = 64'd15;
    end else if ((1'b1 == ap_CS_fsm_state82)) begin
        temp7_address0 = 64'd13;
    end else if ((1'b1 == ap_CS_fsm_state81)) begin
        temp7_address0 = 64'd11;
    end else if ((1'b1 == ap_CS_fsm_state80)) begin
        temp7_address0 = 64'd9;
    end else if ((1'b1 == ap_CS_fsm_state79)) begin
        temp7_address0 = 64'd7;
    end else if ((1'b1 == ap_CS_fsm_state78)) begin
        temp7_address0 = 64'd5;
    end else if ((1'b1 == ap_CS_fsm_state77)) begin
        temp7_address0 = 64'd3;
    end else if ((1'b1 == ap_CS_fsm_state76)) begin
        temp7_address0 = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0;
    end else begin
        temp7_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state84)) begin
        temp7_address1 = 64'd16;
    end else if ((1'b1 == ap_CS_fsm_state83)) begin
        temp7_address1 = 64'd14;
    end else if ((1'b1 == ap_CS_fsm_state82)) begin
        temp7_address1 = 64'd12;
    end else if ((1'b1 == ap_CS_fsm_state81)) begin
        temp7_address1 = 64'd10;
    end else if ((1'b1 == ap_CS_fsm_state80)) begin
        temp7_address1 = 64'd8;
    end else if ((1'b1 == ap_CS_fsm_state79)) begin
        temp7_address1 = 64'd6;
    end else if ((1'b1 == ap_CS_fsm_state78)) begin
        temp7_address1 = 64'd4;
    end else if ((1'b1 == ap_CS_fsm_state77)) begin
        temp7_address1 = 64'd2;
    end else if ((1'b1 == ap_CS_fsm_state76)) begin
        temp7_address1 = 64'd0;
    end else if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1;
    end else begin
        temp7_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state76) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77))) begin
        temp7_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0;
    end else begin
        temp7_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state76) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77))) begin
        temp7_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1;
    end else begin
        temp7_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_we0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0;
    end else begin
        temp7_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        temp7_we1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1;
    end else begin
        temp7_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state20)) begin
        temp_address0 = 64'd17;
    end else if ((1'b1 == ap_CS_fsm_state19)) begin
        temp_address0 = 64'd15;
    end else if ((1'b1 == ap_CS_fsm_state18)) begin
        temp_address0 = 64'd13;
    end else if ((1'b1 == ap_CS_fsm_state17)) begin
        temp_address0 = 64'd11;
    end else if ((1'b1 == ap_CS_fsm_state16)) begin
        temp_address0 = 64'd9;
    end else if ((1'b1 == ap_CS_fsm_state15)) begin
        temp_address0 = 64'd7;
    end else if ((1'b1 == ap_CS_fsm_state14)) begin
        temp_address0 = 64'd5;
    end else if ((1'b1 == ap_CS_fsm_state13)) begin
        temp_address0 = 64'd4;
    end else if ((1'b1 == ap_CS_fsm_state12)) begin
        temp_address0 = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address0;
    end else begin
        temp_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state20)) begin
        temp_address1 = 64'd16;
    end else if ((1'b1 == ap_CS_fsm_state19)) begin
        temp_address1 = 64'd14;
    end else if ((1'b1 == ap_CS_fsm_state18)) begin
        temp_address1 = 64'd12;
    end else if ((1'b1 == ap_CS_fsm_state17)) begin
        temp_address1 = 64'd10;
    end else if ((1'b1 == ap_CS_fsm_state16)) begin
        temp_address1 = 64'd8;
    end else if ((1'b1 == ap_CS_fsm_state15)) begin
        temp_address1 = 64'd6;
    end else if ((1'b1 == ap_CS_fsm_state14)) begin
        temp_address1 = 64'd3;
    end else if ((1'b1 == ap_CS_fsm_state13)) begin
        temp_address1 = 64'd2;
    end else if ((1'b1 == ap_CS_fsm_state12)) begin
        temp_address1 = 64'd0;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_address1;
    end else begin
        temp_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        temp_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce0;
    end else begin
        temp_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        temp_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_ce1;
    end else begin
        temp_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_we0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we0;
    end else begin
        temp_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state11))) begin
        temp_we1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_R_we1;
    end else begin
        temp_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state78))) begin
        uk_admm_V_address0 = 5'd3;
    end else if (((1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state85))) begin
        uk_admm_V_address0 = 5'd17;
    end else if (((1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state84))) begin
        uk_admm_V_address0 = 5'd15;
    end else if (((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state83))) begin
        uk_admm_V_address0 = 5'd13;
    end else if (((1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state82))) begin
        uk_admm_V_address0 = 5'd11;
    end else if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state81))) begin
        uk_admm_V_address0 = 5'd9;
    end else if (((1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state80))) begin
        uk_admm_V_address0 = 5'd7;
    end else if (((1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state79))) begin
        uk_admm_V_address0 = 5'd5;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        uk_admm_V_address0 = 5'd4;
    end else if (((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state77) | ((1'b1 == ap_CS_fsm_state1) & (icmp_ln74_fu_1292_p2 == 1'd0)))) begin
        uk_admm_V_address0 = 5'd1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        uk_admm_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address0;
    end else begin
        uk_admm_V_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state79))) begin
        uk_admm_V_address1 = 5'd4;
    end else if (((1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state85))) begin
        uk_admm_V_address1 = 5'd16;
    end else if (((1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state84))) begin
        uk_admm_V_address1 = 5'd14;
    end else if (((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state83))) begin
        uk_admm_V_address1 = 5'd12;
    end else if (((1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state82))) begin
        uk_admm_V_address1 = 5'd10;
    end else if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state81))) begin
        uk_admm_V_address1 = 5'd8;
    end else if (((1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state80))) begin
        uk_admm_V_address1 = 5'd6;
    end else if ((1'b1 == ap_CS_fsm_state3)) begin
        uk_admm_V_address1 = 5'd3;
    end else if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state78))) begin
        uk_admm_V_address1 = 5'd2;
    end else if (((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state77) | ((1'b1 == ap_CS_fsm_state1) & (icmp_ln74_fu_1292_p2 == 1'd0)))) begin
        uk_admm_V_address1 = 5'd0;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        uk_admm_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_address1;
    end else begin
        uk_admm_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state85) | ((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (icmp_ln74_fu_1292_p2 == 1'd0)))) begin
        uk_admm_V_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        uk_admm_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce0;
    end else begin
        uk_admm_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state85) | ((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (icmp_ln74_fu_1292_p2 == 1'd0)))) begin
        uk_admm_V_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        uk_admm_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_B_ce1;
    end else begin
        uk_admm_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state85)) begin
        uk_admm_V_d0 = select_ln302_59_fu_21376_p3;
    end else if ((1'b1 == ap_CS_fsm_state84)) begin
        uk_admm_V_d0 = select_ln302_57_fu_21238_p3;
    end else if ((1'b1 == ap_CS_fsm_state83)) begin
        uk_admm_V_d0 = select_ln302_55_fu_21100_p3;
    end else if ((1'b1 == ap_CS_fsm_state82)) begin
        uk_admm_V_d0 = select_ln302_53_fu_20962_p3;
    end else if ((1'b1 == ap_CS_fsm_state81)) begin
        uk_admm_V_d0 = select_ln302_51_fu_20824_p3;
    end else if ((1'b1 == ap_CS_fsm_state80)) begin
        uk_admm_V_d0 = select_ln302_49_fu_20686_p3;
    end else if ((1'b1 == ap_CS_fsm_state79)) begin
        uk_admm_V_d0 = select_ln302_47_fu_20548_p3;
    end else if ((1'b1 == ap_CS_fsm_state78)) begin
        uk_admm_V_d0 = select_ln302_45_fu_20410_p3;
    end else if ((1'b1 == ap_CS_fsm_state77)) begin
        uk_admm_V_d0 = select_ln302_43_fu_20272_p3;
    end else begin
        uk_admm_V_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state85)) begin
        uk_admm_V_d1 = select_ln302_58_fu_21307_p3;
    end else if ((1'b1 == ap_CS_fsm_state84)) begin
        uk_admm_V_d1 = select_ln302_56_fu_21169_p3;
    end else if ((1'b1 == ap_CS_fsm_state83)) begin
        uk_admm_V_d1 = select_ln302_54_fu_21031_p3;
    end else if ((1'b1 == ap_CS_fsm_state82)) begin
        uk_admm_V_d1 = select_ln302_52_fu_20893_p3;
    end else if ((1'b1 == ap_CS_fsm_state81)) begin
        uk_admm_V_d1 = select_ln302_50_fu_20755_p3;
    end else if ((1'b1 == ap_CS_fsm_state80)) begin
        uk_admm_V_d1 = select_ln302_48_fu_20617_p3;
    end else if ((1'b1 == ap_CS_fsm_state79)) begin
        uk_admm_V_d1 = select_ln302_46_fu_20479_p3;
    end else if ((1'b1 == ap_CS_fsm_state78)) begin
        uk_admm_V_d1 = select_ln302_44_fu_20341_p3;
    end else if ((1'b1 == ap_CS_fsm_state77)) begin
        uk_admm_V_d1 = select_ln302_42_fu_20203_p3;
    end else begin
        uk_admm_V_d1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state85))) begin
        uk_admm_V_we0 = 1'b1;
    end else begin
        uk_admm_V_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state85))) begin
        uk_admm_V_we1 = 1'b1;
    end else begin
        uk_admm_V_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state36)) begin
        xk_admm_V_0_ap_vld = 1'b1;
    end else begin
        xk_admm_V_0_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state74))) begin
        zk_admm_V_address0 = 5'd17;
    end else if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state73))) begin
        zk_admm_V_address0 = 5'd15;
    end else if (((1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state72))) begin
        zk_admm_V_address0 = 5'd13;
    end else if (((1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state71))) begin
        zk_admm_V_address0 = 5'd11;
    end else if (((1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state70))) begin
        zk_admm_V_address0 = 5'd9;
    end else if (((1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state69))) begin
        zk_admm_V_address0 = 5'd7;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state68))) begin
        zk_admm_V_address0 = 5'd5;
    end else if (((1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state67))) begin
        zk_admm_V_address0 = 5'd3;
    end else if (((1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state66))) begin
        zk_admm_V_address0 = 5'd1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state11))) begin
        zk_admm_V_address0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address0;
    end else begin
        zk_admm_V_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state74))) begin
        zk_admm_V_address1 = 5'd16;
    end else if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state73))) begin
        zk_admm_V_address1 = 5'd14;
    end else if (((1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state72))) begin
        zk_admm_V_address1 = 5'd12;
    end else if (((1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state71))) begin
        zk_admm_V_address1 = 5'd10;
    end else if (((1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state70))) begin
        zk_admm_V_address1 = 5'd8;
    end else if (((1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state69))) begin
        zk_admm_V_address1 = 5'd6;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state68))) begin
        zk_admm_V_address1 = 5'd4;
    end else if (((1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state67))) begin
        zk_admm_V_address1 = 5'd2;
    end else if (((1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state66))) begin
        zk_admm_V_address1 = 5'd0;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state11))) begin
        zk_admm_V_address1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_address1;
    end else begin
        zk_admm_V_address1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        zk_admm_V_ce0 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state11))) begin
        zk_admm_V_ce0 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce0;
    end else begin
        zk_admm_V_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state67))) begin
        zk_admm_V_ce1 = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state11))) begin
        zk_admm_V_ce1 = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_A_ce1;
    end else begin
        zk_admm_V_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        zk_admm_V_d0 = zext_ln50_17_fu_20138_p1;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        zk_admm_V_d0 = zext_ln50_15_fu_19962_p1;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        zk_admm_V_d0 = zext_ln50_13_fu_19786_p1;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        zk_admm_V_d0 = zext_ln50_11_fu_19610_p1;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        zk_admm_V_d0 = zext_ln50_9_fu_19434_p1;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        zk_admm_V_d0 = zext_ln50_7_fu_19258_p1;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        zk_admm_V_d0 = zext_ln50_5_fu_19082_p1;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        zk_admm_V_d0 = zext_ln50_3_fu_18906_p1;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        zk_admm_V_d0 = zext_ln50_1_fu_18730_p1;
    end else begin
        zk_admm_V_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state65)) begin
        zk_admm_V_d1 = zext_ln50_16_fu_20121_p1;
    end else if ((1'b1 == ap_CS_fsm_state64)) begin
        zk_admm_V_d1 = zext_ln50_14_fu_19945_p1;
    end else if ((1'b1 == ap_CS_fsm_state63)) begin
        zk_admm_V_d1 = zext_ln50_12_fu_19769_p1;
    end else if ((1'b1 == ap_CS_fsm_state62)) begin
        zk_admm_V_d1 = zext_ln50_10_fu_19593_p1;
    end else if ((1'b1 == ap_CS_fsm_state61)) begin
        zk_admm_V_d1 = zext_ln50_8_fu_19417_p1;
    end else if ((1'b1 == ap_CS_fsm_state60)) begin
        zk_admm_V_d1 = zext_ln50_6_fu_19241_p1;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        zk_admm_V_d1 = zext_ln50_4_fu_19065_p1;
    end else if ((1'b1 == ap_CS_fsm_state58)) begin
        zk_admm_V_d1 = zext_ln50_2_fu_18889_p1;
    end else if ((1'b1 == ap_CS_fsm_state57)) begin
        zk_admm_V_d1 = zext_ln50_fu_18713_p1;
    end else begin
        zk_admm_V_d1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        zk_admm_V_we0 = 1'b1;
    end else begin
        zk_admm_V_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state65))) begin
        zk_admm_V_we1 = 1'b1;
    end else begin
        zk_admm_V_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (icmp_ln74_fu_1292_p2 == 1'd1))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state18;
        end
        ap_ST_fsm_state18 : begin
            ap_NS_fsm = ap_ST_fsm_state19;
        end
        ap_ST_fsm_state19 : begin
            ap_NS_fsm = ap_ST_fsm_state20;
        end
        ap_ST_fsm_state20 : begin
            ap_NS_fsm = ap_ST_fsm_state21;
        end
        ap_ST_fsm_state21 : begin
            ap_NS_fsm = ap_ST_fsm_state22;
        end
        ap_ST_fsm_state22 : begin
            ap_NS_fsm = ap_ST_fsm_state23;
        end
        ap_ST_fsm_state23 : begin
            ap_NS_fsm = ap_ST_fsm_state24;
        end
        ap_ST_fsm_state24 : begin
            ap_NS_fsm = ap_ST_fsm_state25;
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state26;
        end
        ap_ST_fsm_state26 : begin
            ap_NS_fsm = ap_ST_fsm_state27;
        end
        ap_ST_fsm_state27 : begin
            ap_NS_fsm = ap_ST_fsm_state28;
        end
        ap_ST_fsm_state28 : begin
            ap_NS_fsm = ap_ST_fsm_state29;
        end
        ap_ST_fsm_state29 : begin
            ap_NS_fsm = ap_ST_fsm_state30;
        end
        ap_ST_fsm_state30 : begin
            ap_NS_fsm = ap_ST_fsm_state31;
        end
        ap_ST_fsm_state31 : begin
            ap_NS_fsm = ap_ST_fsm_state32;
        end
        ap_ST_fsm_state32 : begin
            ap_NS_fsm = ap_ST_fsm_state33;
        end
        ap_ST_fsm_state33 : begin
            ap_NS_fsm = ap_ST_fsm_state34;
        end
        ap_ST_fsm_state34 : begin
            ap_NS_fsm = ap_ST_fsm_state35;
        end
        ap_ST_fsm_state35 : begin
            ap_NS_fsm = ap_ST_fsm_state36;
        end
        ap_ST_fsm_state36 : begin
            ap_NS_fsm = ap_ST_fsm_state37;
        end
        ap_ST_fsm_state37 : begin
            ap_NS_fsm = ap_ST_fsm_state38;
        end
        ap_ST_fsm_state38 : begin
            ap_NS_fsm = ap_ST_fsm_state39;
        end
        ap_ST_fsm_state39 : begin
            ap_NS_fsm = ap_ST_fsm_state40;
        end
        ap_ST_fsm_state40 : begin
            ap_NS_fsm = ap_ST_fsm_state41;
        end
        ap_ST_fsm_state41 : begin
            ap_NS_fsm = ap_ST_fsm_state42;
        end
        ap_ST_fsm_state42 : begin
            ap_NS_fsm = ap_ST_fsm_state43;
        end
        ap_ST_fsm_state43 : begin
            ap_NS_fsm = ap_ST_fsm_state44;
        end
        ap_ST_fsm_state44 : begin
            ap_NS_fsm = ap_ST_fsm_state45;
        end
        ap_ST_fsm_state45 : begin
            ap_NS_fsm = ap_ST_fsm_state46;
        end
        ap_ST_fsm_state46 : begin
            ap_NS_fsm = ap_ST_fsm_state47;
        end
        ap_ST_fsm_state47 : begin
            ap_NS_fsm = ap_ST_fsm_state48;
        end
        ap_ST_fsm_state48 : begin
            ap_NS_fsm = ap_ST_fsm_state49;
        end
        ap_ST_fsm_state49 : begin
            ap_NS_fsm = ap_ST_fsm_state50;
        end
        ap_ST_fsm_state50 : begin
            ap_NS_fsm = ap_ST_fsm_state51;
        end
        ap_ST_fsm_state51 : begin
            ap_NS_fsm = ap_ST_fsm_state52;
        end
        ap_ST_fsm_state52 : begin
            ap_NS_fsm = ap_ST_fsm_state53;
        end
        ap_ST_fsm_state53 : begin
            ap_NS_fsm = ap_ST_fsm_state54;
        end
        ap_ST_fsm_state54 : begin
            ap_NS_fsm = ap_ST_fsm_state55;
        end
        ap_ST_fsm_state55 : begin
            ap_NS_fsm = ap_ST_fsm_state56;
        end
        ap_ST_fsm_state56 : begin
            ap_NS_fsm = ap_ST_fsm_state57;
        end
        ap_ST_fsm_state57 : begin
            ap_NS_fsm = ap_ST_fsm_state58;
        end
        ap_ST_fsm_state58 : begin
            ap_NS_fsm = ap_ST_fsm_state59;
        end
        ap_ST_fsm_state59 : begin
            ap_NS_fsm = ap_ST_fsm_state60;
        end
        ap_ST_fsm_state60 : begin
            ap_NS_fsm = ap_ST_fsm_state61;
        end
        ap_ST_fsm_state61 : begin
            ap_NS_fsm = ap_ST_fsm_state62;
        end
        ap_ST_fsm_state62 : begin
            ap_NS_fsm = ap_ST_fsm_state63;
        end
        ap_ST_fsm_state63 : begin
            ap_NS_fsm = ap_ST_fsm_state64;
        end
        ap_ST_fsm_state64 : begin
            ap_NS_fsm = ap_ST_fsm_state65;
        end
        ap_ST_fsm_state65 : begin
            ap_NS_fsm = ap_ST_fsm_state66;
        end
        ap_ST_fsm_state66 : begin
            ap_NS_fsm = ap_ST_fsm_state67;
        end
        ap_ST_fsm_state67 : begin
            ap_NS_fsm = ap_ST_fsm_state68;
        end
        ap_ST_fsm_state68 : begin
            ap_NS_fsm = ap_ST_fsm_state69;
        end
        ap_ST_fsm_state69 : begin
            ap_NS_fsm = ap_ST_fsm_state70;
        end
        ap_ST_fsm_state70 : begin
            ap_NS_fsm = ap_ST_fsm_state71;
        end
        ap_ST_fsm_state71 : begin
            ap_NS_fsm = ap_ST_fsm_state72;
        end
        ap_ST_fsm_state72 : begin
            ap_NS_fsm = ap_ST_fsm_state73;
        end
        ap_ST_fsm_state73 : begin
            ap_NS_fsm = ap_ST_fsm_state74;
        end
        ap_ST_fsm_state74 : begin
            ap_NS_fsm = ap_ST_fsm_state75;
        end
        ap_ST_fsm_state75 : begin
            ap_NS_fsm = ap_ST_fsm_state76;
        end
        ap_ST_fsm_state76 : begin
            ap_NS_fsm = ap_ST_fsm_state77;
        end
        ap_ST_fsm_state77 : begin
            ap_NS_fsm = ap_ST_fsm_state78;
        end
        ap_ST_fsm_state78 : begin
            ap_NS_fsm = ap_ST_fsm_state79;
        end
        ap_ST_fsm_state79 : begin
            ap_NS_fsm = ap_ST_fsm_state80;
        end
        ap_ST_fsm_state80 : begin
            ap_NS_fsm = ap_ST_fsm_state81;
        end
        ap_ST_fsm_state81 : begin
            ap_NS_fsm = ap_ST_fsm_state82;
        end
        ap_ST_fsm_state82 : begin
            ap_NS_fsm = ap_ST_fsm_state83;
        end
        ap_ST_fsm_state83 : begin
            ap_NS_fsm = ap_ST_fsm_state84;
        end
        ap_ST_fsm_state84 : begin
            ap_NS_fsm = ap_ST_fsm_state85;
        end
        ap_ST_fsm_state85 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln1347_10_fu_2939_p2 = ($signed(sext_ln813_56_fu_2935_p1) + $signed(sext_ln813_55_fu_2931_p1));

assign add_ln1347_11_fu_3009_p2 = ($signed(sext_ln813_58_fu_3005_p1) + $signed(sext_ln813_57_fu_3001_p1));

assign add_ln1347_12_fu_3658_p2 = ($signed(sext_ln813_60_fu_3654_p1) + $signed(sext_ln813_59_fu_3650_p1));

assign add_ln1347_13_fu_3728_p2 = ($signed(sext_ln813_62_fu_3724_p1) + $signed(sext_ln813_61_fu_3720_p1));

assign add_ln1347_14_fu_4515_p2 = ($signed(sext_ln813_64_fu_4511_p1) + $signed(sext_ln813_63_fu_4507_p1));

assign add_ln1347_15_fu_4585_p2 = ($signed(sext_ln813_66_fu_4581_p1) + $signed(sext_ln813_65_fu_4577_p1));

assign add_ln1347_16_fu_5150_p2 = ($signed(sext_ln813_68_fu_5146_p1) + $signed(sext_ln813_67_fu_5142_p1));

assign add_ln1347_17_fu_5220_p2 = ($signed(sext_ln813_70_fu_5216_p1) + $signed(sext_ln813_69_fu_5212_p1));

assign add_ln1347_18_fu_2335_p2 = ($signed(sext_ln813_74_fu_2325_p1) + $signed(sext_ln1347_fu_2329_p1));

assign add_ln1347_19_fu_3085_p2 = ($signed(sext_ln813_75_fu_3078_p1) + $signed(sext_ln1347_2_fu_3082_p1));

assign add_ln1347_1_fu_1387_p2 = ($signed(sext_ln813_38_fu_1383_p1) + $signed(sext_ln813_37_fu_1379_p1));

assign add_ln1347_20_fu_3837_p2 = ($signed(sext_ln813_76_fu_3825_p1) + $signed(sext_ln1347_3_fu_3829_p1));

assign add_ln1347_21_fu_4678_p2 = ($signed(sext_ln813_77_fu_4668_p1) + $signed(sext_ln1347_5_fu_4672_p1));

assign add_ln1347_22_fu_5299_p2 = ($signed(sext_ln813_78_fu_5289_p1) + $signed(sext_ln1347_7_fu_5293_p1));

assign add_ln1347_23_fu_5990_p2 = ($signed(sext_ln813_79_fu_5983_p1) + $signed(sext_ln1347_9_fu_5987_p1));

assign add_ln1347_24_fu_6685_p2 = ($signed(sext_ln813_80_fu_6675_p1) + $signed(sext_ln1347_10_fu_6679_p1));

assign add_ln1347_25_fu_7398_p2 = ($signed(sext_ln813_81_fu_7391_p1) + $signed(sext_ln1347_12_fu_7395_p1));

assign add_ln1347_26_fu_8181_p2 = ($signed(sext_ln813_82_fu_8169_p1) + $signed(sext_ln1347_13_fu_8173_p1));

assign add_ln1347_27_fu_8804_p2 = ($signed(sext_ln813_83_fu_8794_p1) + $signed(sext_ln1347_15_fu_8798_p1));

assign add_ln1347_28_fu_9313_p2 = ($signed(sext_ln813_84_fu_9303_p1) + $signed(sext_ln1347_17_fu_9307_p1));

assign add_ln1347_29_fu_9681_p2 = ($signed(sext_ln813_85_fu_9677_p1) + $signed(mul_ln1273_10_reg_22897));

assign add_ln1347_2_fu_1465_p2 = ($signed(sext_ln813_40_fu_1461_p1) + $signed(sext_ln813_39_fu_1457_p1));

assign add_ln1347_30_fu_9992_p2 = ($signed(sext_ln813_86_fu_9988_p1) + $signed(mul_ln1273_11_reg_22952));

assign add_ln1347_31_fu_3319_p2 = ($signed(sext_ln813_87_fu_3309_p1) + $signed(sext_ln1347_19_fu_3313_p1));

assign add_ln1347_32_fu_4087_p2 = ($signed(sext_ln813_88_fu_4080_p1) + $signed(sext_ln1347_21_fu_4084_p1));

assign add_ln1347_33_fu_4945_p2 = ($signed(sext_ln813_89_fu_4933_p1) + $signed(sext_ln1347_22_fu_4937_p1));

assign add_ln1347_34_fu_5636_p2 = ($signed(sext_ln813_90_fu_5629_p1) + $signed(sext_ln1347_24_fu_5633_p1));

assign add_ln1347_35_fu_6247_p2 = ($signed(sext_ln813_91_fu_6237_p1) + $signed(sext_ln1347_25_fu_6241_p1));

assign add_ln1347_36_fu_6915_p2 = ($signed(sext_ln813_92_fu_6908_p1) + $signed(sext_ln1347_27_fu_6912_p1));

assign add_ln1347_37_fu_7639_p2 = ($signed(sext_ln813_93_fu_7627_p1) + $signed(sext_ln1347_28_fu_7631_p1));

assign add_ln1347_38_fu_8444_p2 = ($signed(sext_ln813_94_fu_8440_p1) + $signed(mul_ln1273_18_reg_22922));

assign add_ln1347_39_fu_9124_p2 = ($signed(sext_ln813_95_fu_9120_p1) + $signed(mul_ln1273_19_reg_23023));

assign add_ln1347_3_fu_1617_p2 = ($signed(sext_ln813_42_fu_1613_p1) + $signed(sext_ln813_41_fu_1609_p1));

assign add_ln1347_40_fu_3493_p2 = ($signed(sext_ln813_96_fu_3483_p1) + $signed(sext_ln1347_30_fu_3487_p1));

assign add_ln1347_41_fu_5809_p2 = ($signed(sext_ln813_97_fu_5802_p1) + $signed(sext_ln1347_32_fu_5806_p1));

assign add_ln1347_42_fu_6489_p2 = ($signed(sext_ln813_98_fu_6479_p1) + $signed(sext_ln1347_33_fu_6483_p1));

assign add_ln1347_43_fu_7234_p2 = ($signed(sext_ln813_99_fu_7230_p1) + $signed(grp_fu_21567_p2));

assign add_ln1347_44_fu_7984_p2 = ($signed(sext_ln813_101_fu_7980_p1) + $signed(grp_fu_21582_p2));

assign add_ln1347_45_fu_10924_p2 = ($signed(sext_ln813_104_fu_10914_p1) + $signed(sext_ln1347_35_fu_10918_p1));

assign add_ln1347_46_fu_11599_p2 = ($signed(sext_ln813_105_fu_11589_p1) + $signed(sext_ln1347_37_fu_11593_p1));

assign add_ln1347_47_fu_11154_p2 = ($signed(sext_ln813_106_fu_11144_p1) + $signed(sext_ln1347_39_fu_11148_p1));

assign add_ln1347_48_fu_11795_p2 = ($signed(sext_ln813_107_fu_11785_p1) + $signed(sext_ln1347_41_fu_11789_p1));

assign add_ln1347_49_fu_11403_p2 = ($signed(sext_ln813_108_fu_11391_p1) + $signed(sext_ln1347_43_fu_11395_p1));

assign add_ln1347_4_fu_1535_p2 = ($signed(sext_ln813_44_fu_1531_p1) + $signed(sext_ln813_43_fu_1527_p1));

assign add_ln1347_50_fu_12002_p2 = ($signed(sext_ln813_109_fu_11995_p1) + $signed(sext_ln1347_45_fu_11999_p1));

assign add_ln1347_51_fu_15177_p2 = ($signed(sext_ln813_110_fu_15170_p1) + $signed(sext_ln1347_46_fu_15174_p1));

assign add_ln1347_52_fu_15368_p2 = ($signed(sext_ln813_111_fu_15358_p1) + $signed(sext_ln1347_47_fu_15362_p1));

assign add_ln1347_53_fu_15539_p2 = ($signed(sext_ln813_112_fu_15532_p1) + $signed(sext_ln1347_49_fu_15536_p1));

assign add_ln1347_54_fu_17325_p2 = ($signed(sext_ln813_113_fu_17318_p1) + $signed(sext_ln1347_50_fu_17322_p1));

assign add_ln1347_55_fu_15775_p2 = ($signed(sext_ln813_114_fu_15765_p1) + $signed(sext_ln1347_51_fu_15769_p1));

assign add_ln1347_56_fu_17536_p2 = ($signed(sext_ln813_115_fu_17526_p1) + $signed(sext_ln1347_53_fu_17530_p1));

assign add_ln1347_57_fu_16335_p2 = ($signed(sext_ln813_116_fu_16328_p1) + $signed(sext_ln1347_55_fu_16332_p1));

assign add_ln1347_58_fu_16526_p2 = ($signed(sext_ln813_117_fu_16516_p1) + $signed(sext_ln1347_56_fu_16520_p1));

assign add_ln1347_59_fu_16697_p2 = ($signed(sext_ln813_118_fu_16690_p1) + $signed(sext_ln1347_58_fu_16694_p1));

assign add_ln1347_5_fu_1687_p2 = ($signed(sext_ln813_46_fu_1683_p1) + $signed(sext_ln813_45_fu_1679_p1));

assign add_ln1347_60_fu_18153_p2 = ($signed(sext_ln813_119_fu_18146_p1) + $signed(sext_ln1347_59_fu_18150_p1));

assign add_ln1347_61_fu_16933_p2 = ($signed(sext_ln813_120_fu_16923_p1) + $signed(sext_ln1347_60_fu_16927_p1));

assign add_ln1347_62_fu_18364_p2 = ($signed(sext_ln813_121_fu_18354_p1) + $signed(sext_ln1347_62_fu_18358_p1));

assign add_ln1347_63_fu_18567_p2 = ($signed(sext_ln813_123_fu_18563_p1) + $signed(sext_ln813_122_fu_18559_p1));

assign add_ln1347_64_fu_18638_p2 = ($signed(sext_ln813_125_fu_18634_p1) + $signed(sext_ln813_124_fu_18630_p1));

assign add_ln1347_65_fu_18743_p2 = ($signed(sext_ln813_127_fu_18739_p1) + $signed(sext_ln813_126_fu_18735_p1));

assign add_ln1347_66_fu_18814_p2 = ($signed(sext_ln813_129_fu_18810_p1) + $signed(sext_ln813_128_fu_18806_p1));

assign add_ln1347_67_fu_18919_p2 = ($signed(sext_ln813_131_fu_18915_p1) + $signed(sext_ln813_130_fu_18911_p1));

assign add_ln1347_68_fu_18990_p2 = ($signed(sext_ln813_133_fu_18986_p1) + $signed(sext_ln813_132_fu_18982_p1));

assign add_ln1347_69_fu_19095_p2 = ($signed(sext_ln813_135_fu_19091_p1) + $signed(sext_ln813_134_fu_19087_p1));

assign add_ln1347_6_fu_1845_p2 = ($signed(sext_ln813_48_fu_1841_p1) + $signed(sext_ln813_47_fu_1837_p1));

assign add_ln1347_70_fu_19166_p2 = ($signed(sext_ln813_137_fu_19162_p1) + $signed(sext_ln813_136_fu_19158_p1));

assign add_ln1347_71_fu_19271_p2 = ($signed(sext_ln813_139_fu_19267_p1) + $signed(sext_ln813_138_fu_19263_p1));

assign add_ln1347_72_fu_19342_p2 = ($signed(sext_ln813_141_fu_19338_p1) + $signed(sext_ln813_140_fu_19334_p1));

assign add_ln1347_73_fu_19447_p2 = ($signed(sext_ln813_143_fu_19443_p1) + $signed(sext_ln813_142_fu_19439_p1));

assign add_ln1347_74_fu_19518_p2 = ($signed(sext_ln813_145_fu_19514_p1) + $signed(sext_ln813_144_fu_19510_p1));

assign add_ln1347_75_fu_19623_p2 = ($signed(sext_ln813_147_fu_19619_p1) + $signed(sext_ln813_146_fu_19615_p1));

assign add_ln1347_76_fu_19694_p2 = ($signed(sext_ln813_149_fu_19690_p1) + $signed(sext_ln813_148_fu_19686_p1));

assign add_ln1347_77_fu_19799_p2 = ($signed(sext_ln813_151_fu_19795_p1) + $signed(sext_ln813_150_fu_19791_p1));

assign add_ln1347_78_fu_19870_p2 = ($signed(sext_ln813_153_fu_19866_p1) + $signed(sext_ln813_152_fu_19862_p1));

assign add_ln1347_79_fu_19975_p2 = ($signed(sext_ln813_155_fu_19971_p1) + $signed(sext_ln813_154_fu_19967_p1));

assign add_ln1347_7_fu_1915_p2 = ($signed(sext_ln813_50_fu_1911_p1) + $signed(sext_ln813_49_fu_1907_p1));

assign add_ln1347_80_fu_20046_p2 = ($signed(sext_ln813_157_fu_20042_p1) + $signed(sext_ln813_156_fu_20038_p1));

assign add_ln1347_81_fu_20150_p2 = ($signed(sext_ln813_159_fu_20147_p1) + $signed(sext_ln813_158_fu_20143_p1));

assign add_ln1347_82_fu_20219_p2 = ($signed(sext_ln813_161_fu_20216_p1) + $signed(sext_ln813_160_fu_20212_p1));

assign add_ln1347_83_fu_20288_p2 = ($signed(sext_ln813_163_fu_20285_p1) + $signed(sext_ln813_162_fu_20281_p1));

assign add_ln1347_84_fu_20357_p2 = ($signed(sext_ln813_165_fu_20354_p1) + $signed(sext_ln813_164_fu_20350_p1));

assign add_ln1347_85_fu_20426_p2 = ($signed(sext_ln813_167_fu_20423_p1) + $signed(sext_ln813_166_fu_20419_p1));

assign add_ln1347_86_fu_20495_p2 = ($signed(sext_ln813_169_fu_20492_p1) + $signed(sext_ln813_168_fu_20488_p1));

assign add_ln1347_87_fu_20564_p2 = ($signed(sext_ln813_171_fu_20561_p1) + $signed(sext_ln813_170_fu_20557_p1));

assign add_ln1347_88_fu_20633_p2 = ($signed(sext_ln813_173_fu_20630_p1) + $signed(sext_ln813_172_fu_20626_p1));

assign add_ln1347_89_fu_20702_p2 = ($signed(sext_ln813_175_fu_20699_p1) + $signed(sext_ln813_174_fu_20695_p1));

assign add_ln1347_8_fu_2186_p2 = ($signed(sext_ln813_52_fu_2182_p1) + $signed(sext_ln813_51_fu_2178_p1));

assign add_ln1347_90_fu_20771_p2 = ($signed(sext_ln813_177_fu_20768_p1) + $signed(sext_ln813_176_fu_20764_p1));

assign add_ln1347_91_fu_20840_p2 = ($signed(sext_ln813_179_fu_20837_p1) + $signed(sext_ln813_178_fu_20833_p1));

assign add_ln1347_92_fu_20909_p2 = ($signed(sext_ln813_181_fu_20906_p1) + $signed(sext_ln813_180_fu_20902_p1));

assign add_ln1347_93_fu_20978_p2 = ($signed(sext_ln813_183_fu_20975_p1) + $signed(sext_ln813_182_fu_20971_p1));

assign add_ln1347_94_fu_21047_p2 = ($signed(sext_ln813_185_fu_21044_p1) + $signed(sext_ln813_184_fu_21040_p1));

assign add_ln1347_95_fu_21116_p2 = ($signed(sext_ln813_187_fu_21113_p1) + $signed(sext_ln813_186_fu_21109_p1));

assign add_ln1347_96_fu_21185_p2 = ($signed(sext_ln813_189_fu_21182_p1) + $signed(sext_ln813_188_fu_21178_p1));

assign add_ln1347_97_fu_21254_p2 = ($signed(sext_ln813_191_fu_21251_p1) + $signed(sext_ln813_190_fu_21247_p1));

assign add_ln1347_98_fu_21323_p2 = ($signed(sext_ln813_193_fu_21320_p1) + $signed(sext_ln813_192_fu_21316_p1));

assign add_ln1347_9_fu_2256_p2 = ($signed(sext_ln813_54_fu_2252_p1) + $signed(sext_ln813_53_fu_2248_p1));

assign add_ln1347_fu_1317_p2 = ($signed(sext_ln813_36_fu_1313_p1) + $signed(sext_ln813_fu_1309_p1));

assign add_ln377_10_fu_8845_p2 = (zext_ln377_10_fu_8842_p1 + trunc_ln818_s_fu_8824_p4);

assign add_ln377_11_fu_9354_p2 = (zext_ln377_11_fu_9351_p1 + trunc_ln818_10_fu_9333_p4);

assign add_ln377_12_fu_9715_p2 = (zext_ln377_12_fu_9712_p1 + trunc_ln818_11_fu_9694_p4);

assign add_ln377_13_fu_10026_p2 = (zext_ln377_13_fu_10023_p1 + trunc_ln818_12_fu_10005_p4);

assign add_ln377_14_fu_2586_p2 = (zext_ln377_14_fu_2582_p1 + trunc_ln818_13_fu_2559_p4);

assign add_ln377_15_fu_3368_p2 = (zext_ln377_15_fu_3364_p1 + trunc_ln818_14_fu_3339_p4);

assign add_ln377_16_fu_4127_p2 = (zext_ln377_16_fu_4124_p1 + trunc_ln818_15_fu_4106_p4);

assign add_ln377_17_fu_4986_p2 = (zext_ln377_17_fu_4983_p1 + trunc_ln818_16_fu_4965_p4);

assign add_ln377_18_fu_5676_p2 = (zext_ln377_18_fu_5673_p1 + trunc_ln818_17_fu_5655_p4);

assign add_ln377_19_fu_6288_p2 = (zext_ln377_19_fu_6285_p1 + trunc_ln818_18_fu_6267_p4);

assign add_ln377_1_fu_2376_p2 = (zext_ln377_1_fu_2373_p1 + trunc_ln818_1_fu_2355_p4);

assign add_ln377_20_fu_6955_p2 = (zext_ln377_20_fu_6952_p1 + trunc_ln818_19_fu_6934_p4);

assign add_ln377_21_fu_7689_p2 = (zext_ln377_21_fu_7685_p1 + trunc_ln818_20_fu_7659_p4);

assign add_ln377_22_fu_8478_p2 = (zext_ln377_22_fu_8475_p1 + trunc_ln818_21_fu_8457_p4);

assign add_ln377_23_fu_9158_p2 = (zext_ln377_23_fu_9155_p1 + trunc_ln818_22_fu_9137_p4);

assign add_ln377_24_fu_2779_p2 = (zext_ln377_24_fu_2775_p1 + trunc_ln818_23_fu_2752_p4);

assign add_ln377_25_fu_3542_p2 = (zext_ln377_25_fu_3538_p1 + trunc_ln818_24_fu_3513_p4);

assign add_ln377_26_fu_5857_p2 = (zext_ln377_26_fu_5853_p1 + trunc_ln818_25_fu_5828_p4);

assign add_ln377_27_fu_6530_p2 = (zext_ln377_27_fu_6527_p1 + trunc_ln818_26_fu_6509_p4);

assign add_ln377_28_fu_7276_p2 = (zext_ln377_28_fu_7272_p1 + trunc_ln818_27_fu_7247_p4);

assign add_ln377_29_fu_8026_p2 = (zext_ln377_29_fu_8022_p1 + trunc_ln818_28_fu_7997_p4);

assign add_ln377_2_fu_3125_p2 = (zext_ln377_2_fu_3122_p1 + trunc_ln818_2_fu_3104_p4);

assign add_ln377_30_fu_10404_p2 = ($signed(zext_ln377_30_fu_10400_p1) + $signed(sext_ln818_fu_10382_p1));

assign add_ln377_31_fu_10965_p2 = (zext_ln377_31_fu_10962_p1 + trunc_ln818_30_fu_10944_p4);

assign add_ln377_32_fu_11640_p2 = (zext_ln377_32_fu_11637_p1 + trunc_ln818_31_fu_11619_p4);

assign add_ln377_33_fu_10594_p2 = ($signed(zext_ln377_33_fu_10590_p1) + $signed(sext_ln365_fu_10572_p1));

assign add_ln377_34_fu_11195_p2 = (zext_ln377_34_fu_11192_p1 + trunc_ln818_33_fu_11174_p4);

assign add_ln377_35_fu_11836_p2 = (zext_ln377_35_fu_11833_p1 + trunc_ln818_34_fu_11815_p4);

assign add_ln377_36_fu_10768_p2 = ($signed(zext_ln377_36_fu_10764_p1) + $signed(sext_ln365_1_fu_10746_p1));

assign add_ln377_37_fu_11444_p2 = (zext_ln377_37_fu_11441_p1 + trunc_ln818_36_fu_11423_p4);

assign add_ln377_38_fu_12042_p2 = (zext_ln377_38_fu_12039_p1 + trunc_ln818_37_fu_12021_p4);

assign add_ln377_39_fu_13145_p2 = (zext_ln377_39_fu_13141_p1 + trunc_ln818_38_fu_13118_p4);

assign add_ln377_3_fu_3878_p2 = (zext_ln377_3_fu_3875_p1 + trunc_ln818_3_fu_3857_p4);

assign add_ln377_40_fu_13319_p2 = ($signed(zext_ln377_40_fu_13315_p1) + $signed(sext_ln365_2_fu_13297_p1));

assign add_ln377_41_fu_13489_p2 = (zext_ln377_41_fu_13485_p1 + trunc_ln818_40_fu_13462_p4);

assign add_ln377_42_fu_15225_p2 = (zext_ln377_42_fu_15221_p1 + trunc_ln818_41_fu_15196_p4);

assign add_ln377_43_fu_13679_p2 = ($signed(zext_ln377_43_fu_13675_p1) + $signed(sext_ln365_3_fu_13657_p1));

assign add_ln377_44_fu_15417_p2 = (zext_ln377_44_fu_15413_p1 + trunc_ln818_43_fu_15388_p4);

assign add_ln377_45_fu_13853_p2 = ($signed(zext_ln377_45_fu_13849_p1) + $signed(sext_ln818_1_fu_13831_p1));

assign add_ln377_46_fu_15579_p2 = (zext_ln377_46_fu_15576_p1 + trunc_ln818_45_fu_15558_p4);

assign add_ln377_47_fu_17365_p2 = (zext_ln377_47_fu_17362_p1 + trunc_ln818_46_fu_17344_p4);

assign add_ln377_48_fu_14050_p2 = ($signed(zext_ln377_48_fu_14046_p1) + $signed(sext_ln365_4_fu_14028_p1));

assign add_ln377_49_fu_15816_p2 = (zext_ln377_49_fu_15813_p1 + trunc_ln818_48_fu_15795_p4);

assign add_ln377_4_fu_4719_p2 = (zext_ln377_4_fu_4716_p1 + trunc_ln818_4_fu_4698_p4);

assign add_ln377_50_fu_17577_p2 = (zext_ln377_50_fu_17574_p1 + trunc_ln818_49_fu_17556_p4);

assign add_ln377_51_fu_16011_p2 = (zext_ln377_51_fu_16007_p1 + trunc_ln818_50_fu_15984_p4);

assign add_ln377_52_fu_16185_p2 = ($signed(zext_ln377_52_fu_16181_p1) + $signed(sext_ln365_5_fu_16163_p1));

assign add_ln377_53_fu_14227_p2 = (zext_ln377_53_fu_14223_p1 + trunc_ln818_52_fu_14200_p4);

assign add_ln377_54_fu_16383_p2 = (zext_ln377_54_fu_16379_p1 + trunc_ln818_53_fu_16354_p4);

assign add_ln377_55_fu_14417_p2 = ($signed(zext_ln377_55_fu_14413_p1) + $signed(sext_ln365_6_fu_14395_p1));

assign add_ln377_56_fu_16575_p2 = (zext_ln377_56_fu_16571_p1 + trunc_ln818_55_fu_16546_p4);

assign add_ln377_57_fu_14591_p2 = ($signed(zext_ln377_57_fu_14587_p1) + $signed(sext_ln818_2_fu_14569_p1));

assign add_ln377_58_fu_16737_p2 = (zext_ln377_58_fu_16734_p1 + trunc_ln818_57_fu_16716_p4);

assign add_ln377_59_fu_18193_p2 = (zext_ln377_59_fu_18190_p1 + trunc_ln818_58_fu_18172_p4);

assign add_ln377_5_fu_5340_p2 = (zext_ln377_5_fu_5337_p1 + trunc_ln818_5_fu_5319_p4);

assign add_ln377_60_fu_14788_p2 = ($signed(zext_ln377_60_fu_14784_p1) + $signed(sext_ln365_7_fu_14766_p1));

assign add_ln377_61_fu_16974_p2 = (zext_ln377_61_fu_16971_p1 + trunc_ln818_60_fu_16953_p4);

assign add_ln377_62_fu_18405_p2 = (zext_ln377_62_fu_18402_p1 + trunc_ln818_61_fu_18384_p4);

assign add_ln377_6_fu_6030_p2 = (zext_ln377_6_fu_6027_p1 + trunc_ln818_6_fu_6009_p4);

assign add_ln377_7_fu_6726_p2 = (zext_ln377_7_fu_6723_p1 + trunc_ln818_7_fu_6705_p4);

assign add_ln377_8_fu_7438_p2 = (zext_ln377_8_fu_7435_p1 + trunc_ln818_8_fu_7417_p4);

assign add_ln377_9_fu_8231_p2 = (zext_ln377_9_fu_8227_p1 + trunc_ln818_9_fu_8201_p4);

assign add_ln377_fu_2011_p2 = (zext_ln377_fu_2007_p1 + trunc_ln_fu_1984_p4);

assign add_ln810_10_fu_9319_p2 = ($signed(shl_ln838_s_fu_9296_p3) + $signed(sext_ln1347_18_fu_9310_p1));

assign add_ln810_11_fu_3325_p2 = ($signed(shl_ln838_12_fu_3302_p3) + $signed(sext_ln1347_20_fu_3316_p1));

assign add_ln810_12_fu_4093_p2 = ($signed(shl_ln838_13_fu_4072_p3) + $signed(mul_ln1273_14_reg_22500));

assign add_ln810_13_fu_4951_p2 = ($signed(shl_ln838_14_fu_4925_p3) + $signed(sext_ln1347_23_fu_4941_p1));

assign add_ln810_14_fu_5642_p2 = ($signed(shl_ln838_15_fu_5621_p3) + $signed(mul_ln1273_15_reg_22734));

assign add_ln810_15_fu_6253_p2 = ($signed(shl_ln838_16_fu_6229_p3) + $signed(sext_ln1347_26_fu_6244_p1));

assign add_ln810_16_fu_6921_p2 = ($signed(shl_ln838_17_fu_6900_p3) + $signed(mul_ln1273_17_reg_22824));

assign add_ln810_17_fu_7645_p2 = ($signed(shl_ln838_18_fu_7620_p3) + $signed(sext_ln1347_29_fu_7635_p1));

assign add_ln810_18_fu_3499_p2 = ($signed(shl_ln838_21_fu_3476_p3) + $signed(sext_ln1347_31_fu_3490_p1));

assign add_ln810_19_fu_5815_p2 = ($signed(shl_ln838_22_fu_5795_p3) + $signed(grp_fu_21530_p2));

assign add_ln810_1_fu_3091_p2 = ($signed(shl_ln838_1_fu_3071_p3) + $signed(mul_ln1273_2_reg_22457));

assign add_ln810_20_fu_6495_p2 = ($signed(shl_ln838_23_fu_6471_p3) + $signed(sext_ln1347_34_fu_6486_p1));

assign add_ln810_21_fu_10930_p2 = ($signed(shl_ln838_26_fu_10907_p3) + $signed(sext_ln1347_36_fu_10921_p1));

assign add_ln810_22_fu_11605_p2 = ($signed(shl_ln838_27_fu_11582_p3) + $signed(sext_ln1347_38_fu_11596_p1));

assign add_ln810_23_fu_11160_p2 = ($signed(shl_ln838_28_fu_11136_p3) + $signed(sext_ln1347_40_fu_11151_p1));

assign add_ln810_24_fu_11801_p2 = ($signed(shl_ln838_29_fu_11778_p3) + $signed(sext_ln1347_42_fu_11792_p1));

assign add_ln810_25_fu_11409_p2 = ($signed(shl_ln838_30_fu_11383_p3) + $signed(sext_ln1347_44_fu_11399_p1));

assign add_ln810_26_fu_12008_p2 = ($signed(shl_ln838_31_fu_11987_p3) + $signed(mul_ln1273_32_reg_23202));

assign add_ln810_27_fu_15183_p2 = ($signed(shl_ln838_32_fu_15163_p3) + $signed(grp_fu_21802_p2));

assign add_ln810_28_fu_15374_p2 = ($signed(shl_ln838_33_fu_15350_p3) + $signed(sext_ln1347_48_fu_15365_p1));

assign add_ln810_29_fu_15545_p2 = ($signed(shl_ln838_34_fu_15525_p3) + $signed(mul_ln1273_40_reg_23500));

assign add_ln810_2_fu_3843_p2 = ($signed(shl_ln838_2_fu_3818_p3) + $signed(sext_ln1347_4_fu_3833_p1));

assign add_ln810_30_fu_17331_p2 = ($signed(shl_ln838_35_fu_17311_p3) + $signed(mul_ln1273_41_reg_23676));

assign add_ln810_31_fu_15781_p2 = ($signed(shl_ln838_36_fu_15757_p3) + $signed(sext_ln1347_52_fu_15772_p1));

assign add_ln810_32_fu_17542_p2 = ($signed(shl_ln838_37_fu_17519_p3) + $signed(sext_ln1347_54_fu_17533_p1));

assign add_ln810_33_fu_16341_p2 = ($signed(shl_ln838_38_fu_16321_p3) + $signed(grp_fu_21855_p2));

assign add_ln810_34_fu_16532_p2 = ($signed(shl_ln838_39_fu_16508_p3) + $signed(sext_ln1347_57_fu_16523_p1));

assign add_ln810_35_fu_16703_p2 = ($signed(shl_ln838_40_fu_16683_p3) + $signed(mul_ln1273_52_reg_23562));

assign add_ln810_36_fu_18159_p2 = ($signed(shl_ln838_41_fu_18139_p3) + $signed(mul_ln1273_53_reg_23810));

assign add_ln810_37_fu_16939_p2 = ($signed(shl_ln838_42_fu_16915_p3) + $signed(sext_ln1347_61_fu_16930_p1));

assign add_ln810_38_fu_18370_p2 = ($signed(shl_ln838_43_fu_18347_p3) + $signed(sext_ln1347_63_fu_18361_p1));

assign add_ln810_3_fu_4684_p2 = ($signed(shl_ln838_3_fu_4660_p3) + $signed(sext_ln1347_6_fu_4675_p1));

assign add_ln810_4_fu_5305_p2 = ($signed(shl_ln838_4_fu_5282_p3) + $signed(sext_ln1347_8_fu_5296_p1));

assign add_ln810_5_fu_5996_p2 = ($signed(shl_ln838_5_fu_5976_p3) + $signed(mul_ln1273_5_reg_22646));

assign add_ln810_6_fu_6691_p2 = ($signed(shl_ln838_6_fu_6668_p3) + $signed(sext_ln1347_11_fu_6682_p1));

assign add_ln810_7_fu_7404_p2 = ($signed(shl_ln838_7_fu_7384_p3) + $signed(mul_ln1273_7_reg_22703));

assign add_ln810_8_fu_8187_p2 = ($signed(shl_ln838_8_fu_8162_p3) + $signed(sext_ln1347_14_fu_8177_p1));

assign add_ln810_9_fu_8810_p2 = ($signed(shl_ln838_9_fu_8786_p3) + $signed(sext_ln1347_16_fu_8801_p1));

assign add_ln810_fu_2341_p2 = ($signed(shl_ln_fu_2318_p3) + $signed(sext_ln1347_1_fu_2332_p1));

assign add_ln813_10_fu_2953_p1 = temp_q1;

assign add_ln813_10_fu_2953_p2 = ($signed(reg_1240) + $signed(add_ln813_10_fu_2953_p1));

assign add_ln813_11_fu_3023_p1 = temp_q0;

assign add_ln813_11_fu_3023_p2 = ($signed(reg_1244) + $signed(add_ln813_11_fu_3023_p1));

assign add_ln813_12_fu_3672_p1 = temp_q1;

assign add_ln813_12_fu_3672_p2 = ($signed(reg_1248) + $signed(add_ln813_12_fu_3672_p1));

assign add_ln813_13_fu_3742_p1 = temp_q0;

assign add_ln813_13_fu_3742_p2 = ($signed(reg_1252) + $signed(add_ln813_13_fu_3742_p1));

assign add_ln813_14_fu_4529_p1 = temp_q1;

assign add_ln813_14_fu_4529_p2 = ($signed(reg_1256) + $signed(add_ln813_14_fu_4529_p1));

assign add_ln813_15_fu_4599_p1 = temp_q0;

assign add_ln813_15_fu_4599_p2 = ($signed(reg_1260) + $signed(add_ln813_15_fu_4599_p1));

assign add_ln813_16_fu_5164_p1 = temp_q1;

assign add_ln813_16_fu_5164_p2 = ($signed(reg_1264) + $signed(add_ln813_16_fu_5164_p1));

assign add_ln813_17_fu_5234_p1 = temp_q0;

assign add_ln813_17_fu_5234_p2 = ($signed(reg_1268) + $signed(add_ln813_17_fu_5234_p1));

assign add_ln813_18_fu_18581_p0 = Hxk_V_q1;

assign add_ln813_18_fu_18581_p2 = ($signed(add_ln813_18_fu_18581_p0) + $signed(reg_1200));

assign add_ln813_19_fu_18652_p0 = Hxk_V_q0;

assign add_ln813_19_fu_18652_p2 = ($signed(add_ln813_19_fu_18652_p0) + $signed(reg_1204));

assign add_ln813_1_fu_1401_p1 = temp_q0;

assign add_ln813_1_fu_1401_p2 = ($signed(reg_1204) + $signed(add_ln813_1_fu_1401_p1));

assign add_ln813_20_fu_18757_p0 = Hxk_V_q1;

assign add_ln813_20_fu_18757_p2 = ($signed(add_ln813_20_fu_18757_p0) + $signed(reg_1208));

assign add_ln813_21_fu_18828_p0 = Hxk_V_q0;

assign add_ln813_21_fu_18828_p2 = ($signed(add_ln813_21_fu_18828_p0) + $signed(reg_1212));

assign add_ln813_22_fu_18933_p0 = Hxk_V_q1;

assign add_ln813_22_fu_18933_p2 = ($signed(add_ln813_22_fu_18933_p0) + $signed(reg_1216));

assign add_ln813_23_fu_19004_p0 = Hxk_V_q0;

assign add_ln813_23_fu_19004_p2 = ($signed(add_ln813_23_fu_19004_p0) + $signed(reg_1220));

assign add_ln813_24_fu_19109_p0 = Hxk_V_q1;

assign add_ln813_24_fu_19109_p2 = ($signed(add_ln813_24_fu_19109_p0) + $signed(reg_1224));

assign add_ln813_25_fu_19180_p0 = Hxk_V_q0;

assign add_ln813_25_fu_19180_p2 = ($signed(add_ln813_25_fu_19180_p0) + $signed(reg_1228));

assign add_ln813_26_fu_19285_p0 = Hxk_V_q1;

assign add_ln813_26_fu_19285_p2 = ($signed(add_ln813_26_fu_19285_p0) + $signed(reg_1232));

assign add_ln813_27_fu_19356_p0 = Hxk_V_q0;

assign add_ln813_27_fu_19356_p2 = ($signed(add_ln813_27_fu_19356_p0) + $signed(reg_1236));

assign add_ln813_28_fu_19461_p0 = Hxk_V_q1;

assign add_ln813_28_fu_19461_p2 = ($signed(add_ln813_28_fu_19461_p0) + $signed(reg_1240));

assign add_ln813_29_fu_19532_p0 = Hxk_V_q0;

assign add_ln813_29_fu_19532_p2 = ($signed(add_ln813_29_fu_19532_p0) + $signed(reg_1244));

assign add_ln813_2_fu_1479_p1 = temp_q1;

assign add_ln813_2_fu_1479_p2 = ($signed(reg_1208) + $signed(add_ln813_2_fu_1479_p1));

assign add_ln813_30_fu_19637_p0 = Hxk_V_q1;

assign add_ln813_30_fu_19637_p2 = ($signed(add_ln813_30_fu_19637_p0) + $signed(reg_1248));

assign add_ln813_31_fu_19708_p0 = Hxk_V_q0;

assign add_ln813_31_fu_19708_p2 = ($signed(add_ln813_31_fu_19708_p0) + $signed(reg_1252));

assign add_ln813_32_fu_19813_p0 = Hxk_V_q1;

assign add_ln813_32_fu_19813_p2 = ($signed(add_ln813_32_fu_19813_p0) + $signed(reg_1256));

assign add_ln813_33_fu_19884_p0 = Hxk_V_q0;

assign add_ln813_33_fu_19884_p2 = ($signed(add_ln813_33_fu_19884_p0) + $signed(reg_1260));

assign add_ln813_34_fu_19989_p0 = Hxk_V_q1;

assign add_ln813_34_fu_19989_p2 = ($signed(add_ln813_34_fu_19989_p0) + $signed(reg_1264));

assign add_ln813_35_fu_20060_p0 = Hxk_V_q0;

assign add_ln813_35_fu_20060_p2 = ($signed(add_ln813_35_fu_20060_p0) + $signed(reg_1268));

assign add_ln813_36_fu_20164_p1 = temp7_q1;

assign add_ln813_36_fu_20164_p2 = ($signed(zk_admm_V_load_reg_23882) + $signed(add_ln813_36_fu_20164_p1));

assign add_ln813_37_fu_20233_p1 = temp7_q0;

assign add_ln813_37_fu_20233_p2 = ($signed(zk_admm_V_load_1_reg_23888) + $signed(add_ln813_37_fu_20233_p1));

assign add_ln813_38_fu_20302_p1 = temp7_q1;

assign add_ln813_38_fu_20302_p2 = ($signed(zk_admm_V_load_2_reg_23894) + $signed(add_ln813_38_fu_20302_p1));

assign add_ln813_39_fu_20371_p1 = temp7_q0;

assign add_ln813_39_fu_20371_p2 = ($signed(zk_admm_V_load_3_reg_23900) + $signed(add_ln813_39_fu_20371_p1));

assign add_ln813_3_fu_1631_p1 = temp_q1;

assign add_ln813_3_fu_1631_p2 = ($signed(reg_1216) + $signed(add_ln813_3_fu_1631_p1));

assign add_ln813_40_fu_20440_p1 = temp7_q1;

assign add_ln813_40_fu_20440_p2 = ($signed(zk_admm_V_load_4_reg_23906) + $signed(add_ln813_40_fu_20440_p1));

assign add_ln813_41_fu_20509_p1 = temp7_q0;

assign add_ln813_41_fu_20509_p2 = ($signed(zk_admm_V_load_5_reg_23912) + $signed(add_ln813_41_fu_20509_p1));

assign add_ln813_42_fu_20578_p1 = temp7_q1;

assign add_ln813_42_fu_20578_p2 = ($signed(zk_admm_V_load_6_reg_23918) + $signed(add_ln813_42_fu_20578_p1));

assign add_ln813_43_fu_20647_p1 = temp7_q0;

assign add_ln813_43_fu_20647_p2 = ($signed(zk_admm_V_load_7_reg_23924) + $signed(add_ln813_43_fu_20647_p1));

assign add_ln813_44_fu_20716_p1 = temp7_q1;

assign add_ln813_44_fu_20716_p2 = ($signed(zk_admm_V_load_8_reg_23930) + $signed(add_ln813_44_fu_20716_p1));

assign add_ln813_45_fu_20785_p1 = temp7_q0;

assign add_ln813_45_fu_20785_p2 = ($signed(zk_admm_V_load_9_reg_23936) + $signed(add_ln813_45_fu_20785_p1));

assign add_ln813_46_fu_20854_p1 = temp7_q1;

assign add_ln813_46_fu_20854_p2 = ($signed(zk_admm_V_load_10_reg_23942) + $signed(add_ln813_46_fu_20854_p1));

assign add_ln813_47_fu_20923_p1 = temp7_q0;

assign add_ln813_47_fu_20923_p2 = ($signed(zk_admm_V_load_11_reg_23948) + $signed(add_ln813_47_fu_20923_p1));

assign add_ln813_48_fu_20992_p1 = temp7_q1;

assign add_ln813_48_fu_20992_p2 = ($signed(zk_admm_V_load_12_reg_23954) + $signed(add_ln813_48_fu_20992_p1));

assign add_ln813_49_fu_21061_p1 = temp7_q0;

assign add_ln813_49_fu_21061_p2 = ($signed(zk_admm_V_load_13_reg_23960) + $signed(add_ln813_49_fu_21061_p1));

assign add_ln813_4_fu_1549_p1 = temp_q0;

assign add_ln813_4_fu_1549_p2 = ($signed(reg_1212) + $signed(add_ln813_4_fu_1549_p1));

assign add_ln813_50_fu_21130_p1 = temp7_q1;

assign add_ln813_50_fu_21130_p2 = ($signed(zk_admm_V_load_14_reg_23966) + $signed(add_ln813_50_fu_21130_p1));

assign add_ln813_51_fu_21199_p1 = temp7_q0;

assign add_ln813_51_fu_21199_p2 = ($signed(zk_admm_V_load_15_reg_23972) + $signed(add_ln813_51_fu_21199_p1));

assign add_ln813_52_fu_21268_p1 = temp7_q1;

assign add_ln813_52_fu_21268_p2 = ($signed(zk_admm_V_load_16_reg_23978) + $signed(add_ln813_52_fu_21268_p1));

assign add_ln813_53_fu_21337_p1 = temp7_q0;

assign add_ln813_53_fu_21337_p2 = ($signed(zk_admm_V_load_17_reg_23984) + $signed(add_ln813_53_fu_21337_p1));

assign add_ln813_5_fu_1701_p1 = temp_q0;

assign add_ln813_5_fu_1701_p2 = ($signed(reg_1220) + $signed(add_ln813_5_fu_1701_p1));

assign add_ln813_6_fu_1859_p1 = temp_q1;

assign add_ln813_6_fu_1859_p2 = ($signed(reg_1224) + $signed(add_ln813_6_fu_1859_p1));

assign add_ln813_7_fu_1929_p1 = temp_q0;

assign add_ln813_7_fu_1929_p2 = ($signed(reg_1228) + $signed(add_ln813_7_fu_1929_p1));

assign add_ln813_8_fu_2200_p1 = temp_q1;

assign add_ln813_8_fu_2200_p2 = ($signed(reg_1232) + $signed(add_ln813_8_fu_2200_p1));

assign add_ln813_9_fu_2270_p1 = temp_q0;

assign add_ln813_9_fu_2270_p2 = ($signed(reg_1236) + $signed(add_ln813_9_fu_2270_p1));

assign add_ln813_fu_1331_p1 = temp_q1;

assign add_ln813_fu_1331_p2 = ($signed(reg_1200) + $signed(add_ln813_fu_1331_p1));

assign and_ln378_10_fu_8865_p2 = (xor_ln896_20_fu_8859_p2 & tmp_132_fu_8834_p3);

assign and_ln378_11_fu_9374_p2 = (xor_ln896_22_fu_9368_p2 & tmp_138_fu_9343_p3);

assign and_ln378_12_fu_9735_p2 = (xor_ln896_24_fu_9729_p2 & tmp_144_fu_9704_p3);

assign and_ln378_13_fu_10046_p2 = (xor_ln896_28_fu_10040_p2 & tmp_154_fu_10015_p3);

assign and_ln378_14_fu_2606_p2 = (xor_ln896_32_fu_2600_p2 & tmp_164_fu_2568_p3);

assign and_ln378_15_fu_4034_p2 = (xor_ln896_34_reg_22574 & tmp_170_reg_22564);

assign and_ln378_16_fu_4147_p2 = (xor_ln896_36_fu_4141_p2 & tmp_176_fu_4116_p3);

assign and_ln378_17_fu_5006_p2 = (xor_ln896_38_fu_5000_p2 & tmp_182_fu_4975_p3);

assign and_ln378_18_fu_6191_p2 = (xor_ln896_42_reg_22803 & tmp_192_reg_22793);

assign and_ln378_19_fu_6308_p2 = (xor_ln896_44_fu_6302_p2 & tmp_198_fu_6277_p3);

assign and_ln378_1_fu_2396_p2 = (xor_ln896_2_fu_2390_p2 & tmp_78_fu_2365_p3);

assign and_ln378_20_fu_6975_p2 = (xor_ln896_46_fu_6969_p2 & tmp_204_fu_6944_p3);

assign and_ln378_21_fu_7709_p2 = (xor_ln896_48_fu_7703_p2 & tmp_210_fu_7669_p3);

assign and_ln378_22_fu_8498_p2 = (xor_ln896_51_fu_8492_p2 & tmp_218_fu_8467_p3);

assign and_ln378_23_fu_9178_p2 = (xor_ln896_55_fu_9172_p2 & tmp_228_fu_9147_p3);

assign and_ln378_24_fu_2799_p2 = (xor_ln896_58_fu_2793_p2 & tmp_236_fu_2761_p3);

assign and_ln378_25_fu_4269_p2 = (xor_ln896_60_reg_22610 & tmp_242_reg_22600);

assign and_ln378_26_fu_6433_p2 = (xor_ln896_66_reg_22855 & tmp_256_reg_22845);

assign and_ln378_27_fu_6550_p2 = (xor_ln896_68_fu_6544_p2 & tmp_262_fu_6519_p3);

assign and_ln378_28_fu_7834_p2 = (xor_ln896_72_reg_22982 & tmp_272_reg_22972);

assign and_ln378_29_fu_8616_p2 = (xor_ln896_76_reg_23048 & tmp_282_reg_23038);

assign and_ln378_2_fu_3145_p2 = (xor_ln896_4_fu_3139_p2 & tmp_84_fu_3114_p3);

assign and_ln378_30_fu_10424_p2 = (xor_ln896_78_fu_10418_p2 & tmp_294_fu_10386_p3);

assign and_ln378_31_fu_10985_p2 = (xor_ln896_80_fu_10979_p2 & tmp_300_fu_10954_p3);

assign and_ln378_32_fu_11660_p2 = (xor_ln896_82_fu_11654_p2 & tmp_306_fu_11629_p3);

assign and_ln378_33_fu_10614_p2 = (xor_ln896_84_fu_10608_p2 & tmp_312_fu_10576_p3);

assign and_ln378_34_fu_11215_p2 = (xor_ln896_86_fu_11209_p2 & tmp_318_fu_11184_p3);

assign and_ln378_35_fu_11856_p2 = (xor_ln896_88_fu_11850_p2 & tmp_324_fu_11825_p3);

assign and_ln378_36_fu_10788_p2 = (xor_ln896_90_fu_10782_p2 & tmp_330_fu_10750_p3);

assign and_ln378_37_fu_11464_p2 = (xor_ln896_92_fu_11458_p2 & tmp_336_fu_11433_p3);

assign and_ln378_38_fu_12062_p2 = (xor_ln896_94_fu_12056_p2 & tmp_342_fu_12031_p3);

assign and_ln378_39_fu_13165_p2 = (xor_ln896_96_fu_13159_p2 & tmp_348_fu_13127_p3);

assign and_ln378_3_fu_3898_p2 = (xor_ln896_6_fu_3892_p2 & tmp_90_fu_3867_p3);

assign and_ln378_40_fu_13339_p2 = (xor_ln896_100_fu_13333_p2 & tmp_358_fu_13301_p3);

assign and_ln378_41_fu_13509_p2 = (xor_ln896_104_fu_13503_p2 & tmp_368_fu_13471_p3);

assign and_ln378_42_fu_17135_p2 = (xor_ln896_106_reg_23619 & tmp_374_reg_23609);

assign and_ln378_43_fu_13699_p2 = (xor_ln896_109_fu_13693_p2 & tmp_382_fu_13661_p3);

assign and_ln378_44_fu_17223_p2 = (xor_ln896_111_reg_23655 & tmp_388_reg_23645);

assign and_ln378_45_fu_13873_p2 = (xor_ln896_114_fu_13867_p2 & tmp_396_fu_13835_p3);

assign and_ln378_46_fu_15599_p2 = (xor_ln896_116_fu_15593_p2 & tmp_402_fu_15568_p3);

assign and_ln378_47_fu_17385_p2 = (xor_ln896_118_fu_17379_p2 & tmp_408_fu_17354_p3);

assign and_ln378_48_fu_14070_p2 = (xor_ln896_120_fu_14064_p2 & tmp_414_fu_14032_p3);

assign and_ln378_49_fu_15836_p2 = (xor_ln896_122_fu_15830_p2 & tmp_420_fu_15805_p3);

assign and_ln378_4_fu_4739_p2 = (xor_ln896_8_fu_4733_p2 & tmp_96_fu_4708_p3);

assign and_ln378_50_fu_17597_p2 = (xor_ln896_124_fu_17591_p2 & tmp_426_fu_17566_p3);

assign and_ln378_51_fu_16031_p2 = (xor_ln896_126_fu_16025_p2 & tmp_432_fu_15993_p3);

assign and_ln378_52_fu_16205_p2 = (xor_ln896_130_fu_16199_p2 & tmp_442_fu_16167_p3);

assign and_ln378_53_fu_14247_p2 = (xor_ln896_134_fu_14241_p2 & tmp_452_fu_14209_p3);

assign and_ln378_54_fu_17963_p2 = (xor_ln896_136_reg_23753 & tmp_458_reg_23743);

assign and_ln378_55_fu_14437_p2 = (xor_ln896_139_fu_14431_p2 & tmp_466_fu_14399_p3);

assign and_ln378_56_fu_18051_p2 = (xor_ln896_141_reg_23789 & tmp_472_reg_23779);

assign and_ln378_57_fu_14611_p2 = (xor_ln896_144_fu_14605_p2 & tmp_480_fu_14573_p3);

assign and_ln378_58_fu_16757_p2 = (xor_ln896_146_fu_16751_p2 & tmp_486_fu_16726_p3);

assign and_ln378_59_fu_18213_p2 = (xor_ln896_148_fu_18207_p2 & tmp_492_fu_18182_p3);

assign and_ln378_5_fu_5360_p2 = (xor_ln896_10_fu_5354_p2 & tmp_102_fu_5329_p3);

assign and_ln378_60_fu_14808_p2 = (xor_ln896_150_fu_14802_p2 & tmp_498_fu_14770_p3);

assign and_ln378_61_fu_16994_p2 = (xor_ln896_152_fu_16988_p2 & tmp_504_fu_16963_p3);

assign and_ln378_62_fu_18425_p2 = (xor_ln896_154_fu_18419_p2 & tmp_510_fu_18394_p3);

assign and_ln378_6_fu_6050_p2 = (xor_ln896_12_fu_6044_p2 & tmp_108_fu_6019_p3);

assign and_ln378_7_fu_6746_p2 = (xor_ln896_14_fu_6740_p2 & tmp_114_fu_6715_p3);

assign and_ln378_8_fu_7458_p2 = (xor_ln896_16_fu_7452_p2 & tmp_120_fu_7427_p3);

assign and_ln378_9_fu_8251_p2 = (xor_ln896_18_fu_8245_p2 & tmp_126_fu_8211_p3);

assign and_ln378_fu_2031_p2 = (xor_ln896_fu_2025_p2 & tmp_72_fu_1993_p3);

assign and_ln890_10_fu_8917_p2 = (tmp_135_fu_8871_p3 & or_ln890_10_fu_8911_p2);

assign and_ln890_11_fu_9426_p2 = (tmp_141_fu_9380_p3 & or_ln890_11_fu_9420_p2);

assign and_ln890_12_fu_9787_p2 = (tmp_147_fu_9741_p3 & or_ln890_12_fu_9781_p2);

assign and_ln890_13_fu_10098_p2 = (tmp_157_fu_10052_p3 & or_ln890_13_fu_10092_p2);

assign and_ln890_14_fu_2656_p2 = (tmp_167_fu_2612_p3 & or_ln890_14_fu_2650_p2);

assign and_ln890_15_fu_3434_p2 = (tmp_173_fu_3388_p3 & or_ln890_15_fu_3428_p2);

assign and_ln890_16_fu_4199_p2 = (tmp_179_fu_4153_p3 & or_ln890_16_fu_4193_p2);

assign and_ln890_17_fu_5058_p2 = (tmp_185_fu_5012_p3 & or_ln890_17_fu_5052_p2);

assign and_ln890_18_fu_5742_p2 = (tmp_195_fu_5696_p3 & or_ln890_18_fu_5736_p2);

assign and_ln890_19_fu_6360_p2 = (tmp_201_fu_6314_p3 & or_ln890_19_fu_6354_p2);

assign and_ln890_1_fu_2448_p2 = (tmp_81_fu_2402_p3 & or_ln890_1_fu_2442_p2);

assign and_ln890_20_fu_7027_p2 = (tmp_207_fu_6981_p3 & or_ln890_20_fu_7021_p2);

assign and_ln890_21_fu_7761_p2 = (tmp_213_fu_7715_p3 & or_ln890_21_fu_7755_p2);

assign and_ln890_22_fu_8550_p2 = (tmp_221_fu_8504_p3 & or_ln890_22_fu_8544_p2);

assign and_ln890_23_fu_9230_p2 = (tmp_231_fu_9184_p3 & or_ln890_23_fu_9224_p2);

assign and_ln890_24_fu_2849_p2 = (tmp_239_fu_2805_p3 & or_ln890_24_fu_2843_p2);

assign and_ln890_25_fu_3608_p2 = (tmp_245_fu_3562_p3 & or_ln890_25_fu_3602_p2);

assign and_ln890_26_fu_5923_p2 = (tmp_259_fu_5877_p3 & or_ln890_26_fu_5917_p2);

assign and_ln890_27_fu_6602_p2 = (tmp_265_fu_6556_p3 & or_ln890_27_fu_6596_p2);

assign and_ln890_28_fu_7342_p2 = (tmp_275_fu_7296_p3 & or_ln890_28_fu_7336_p2);

assign and_ln890_29_fu_8092_p2 = (tmp_285_fu_8046_p3 & or_ln890_29_fu_8086_p2);

assign and_ln890_2_fu_3197_p2 = (tmp_87_fu_3151_p3 & or_ln890_2_fu_3191_p2);

assign and_ln890_30_fu_10474_p2 = (tmp_297_fu_10430_p3 & or_ln890_30_fu_10468_p2);

assign and_ln890_31_fu_11037_p2 = (tmp_303_fu_10991_p3 & or_ln890_31_fu_11031_p2);

assign and_ln890_32_fu_11712_p2 = (tmp_309_fu_11666_p3 & or_ln890_32_fu_11706_p2);

assign and_ln890_33_fu_10664_p2 = (tmp_315_fu_10620_p3 & or_ln890_33_fu_10658_p2);

assign and_ln890_34_fu_11267_p2 = (tmp_321_fu_11221_p3 & or_ln890_34_fu_11261_p2);

assign and_ln890_35_fu_11908_p2 = (tmp_327_fu_11862_p3 & or_ln890_35_fu_11902_p2);

assign and_ln890_36_fu_10838_p2 = (tmp_333_fu_10794_p3 & or_ln890_36_fu_10832_p2);

assign and_ln890_37_fu_11516_p2 = (tmp_339_fu_11470_p3 & or_ln890_37_fu_11510_p2);

assign and_ln890_38_fu_12114_p2 = (tmp_345_fu_12068_p3 & or_ln890_38_fu_12108_p2);

assign and_ln890_39_fu_13215_p2 = (tmp_351_fu_13171_p3 & or_ln890_39_fu_13209_p2);

assign and_ln890_3_fu_3950_p2 = (tmp_93_fu_3904_p3 & or_ln890_3_fu_3944_p2);

assign and_ln890_40_fu_13389_p2 = (tmp_361_fu_13345_p3 & or_ln890_40_fu_13383_p2);

assign and_ln890_41_fu_13559_p2 = (tmp_371_fu_13515_p3 & or_ln890_41_fu_13553_p2);

assign and_ln890_42_fu_15291_p2 = (tmp_377_fu_15245_p3 & or_ln890_42_fu_15285_p2);

assign and_ln890_43_fu_13749_p2 = (tmp_385_fu_13705_p3 & or_ln890_43_fu_13743_p2);

assign and_ln890_44_fu_15483_p2 = (tmp_391_fu_15437_p3 & or_ln890_44_fu_15477_p2);

assign and_ln890_45_fu_13923_p2 = (tmp_399_fu_13879_p3 & or_ln890_45_fu_13917_p2);

assign and_ln890_46_fu_15651_p2 = (tmp_405_fu_15605_p3 & or_ln890_46_fu_15645_p2);

assign and_ln890_47_fu_17437_p2 = (tmp_411_fu_17391_p3 & or_ln890_47_fu_17431_p2);

assign and_ln890_48_fu_14120_p2 = (tmp_417_fu_14076_p3 & or_ln890_48_fu_14114_p2);

assign and_ln890_49_fu_15888_p2 = (tmp_423_fu_15842_p3 & or_ln890_49_fu_15882_p2);

assign and_ln890_4_fu_4791_p2 = (tmp_99_fu_4745_p3 & or_ln890_4_fu_4785_p2);

assign and_ln890_50_fu_17649_p2 = (tmp_429_fu_17603_p3 & or_ln890_50_fu_17643_p2);

assign and_ln890_51_fu_16081_p2 = (tmp_435_fu_16037_p3 & or_ln890_51_fu_16075_p2);

assign and_ln890_52_fu_16255_p2 = (tmp_445_fu_16211_p3 & or_ln890_52_fu_16249_p2);

assign and_ln890_53_fu_14297_p2 = (tmp_455_fu_14253_p3 & or_ln890_53_fu_14291_p2);

assign and_ln890_54_fu_16449_p2 = (tmp_461_fu_16403_p3 & or_ln890_54_fu_16443_p2);

assign and_ln890_55_fu_14487_p2 = (tmp_469_fu_14443_p3 & or_ln890_55_fu_14481_p2);

assign and_ln890_56_fu_16641_p2 = (tmp_475_fu_16595_p3 & or_ln890_56_fu_16635_p2);

assign and_ln890_57_fu_14661_p2 = (tmp_483_fu_14617_p3 & or_ln890_57_fu_14655_p2);

assign and_ln890_58_fu_16809_p2 = (tmp_489_fu_16763_p3 & or_ln890_58_fu_16803_p2);

assign and_ln890_59_fu_18265_p2 = (tmp_495_fu_18219_p3 & or_ln890_59_fu_18259_p2);

assign and_ln890_5_fu_5412_p2 = (tmp_105_fu_5366_p3 & or_ln890_5_fu_5406_p2);

assign and_ln890_60_fu_14858_p2 = (tmp_501_fu_14814_p3 & or_ln890_60_fu_14852_p2);

assign and_ln890_61_fu_17046_p2 = (tmp_507_fu_17000_p3 & or_ln890_61_fu_17040_p2);

assign and_ln890_62_fu_18477_p2 = (tmp_513_fu_18431_p3 & or_ln890_62_fu_18471_p2);

assign and_ln890_6_fu_6102_p2 = (tmp_111_fu_6056_p3 & or_ln890_6_fu_6096_p2);

assign and_ln890_7_fu_6798_p2 = (tmp_117_fu_6752_p3 & or_ln890_7_fu_6792_p2);

assign and_ln890_8_fu_7510_p2 = (tmp_123_fu_7464_p3 & or_ln890_8_fu_7504_p2);

assign and_ln890_9_fu_8303_p2 = (tmp_129_fu_8257_p3 & or_ln890_9_fu_8297_p2);

assign and_ln890_fu_2081_p2 = (tmp_75_fu_2037_p3 & or_ln890_fu_2075_p2);

assign and_ln891_10_fu_8923_p2 = (tmp_135_fu_8871_p3 & and_ln378_10_fu_8865_p2);

assign and_ln891_11_fu_9432_p2 = (tmp_141_fu_9380_p3 & and_ln378_11_fu_9374_p2);

assign and_ln891_12_fu_9793_p2 = (tmp_147_fu_9741_p3 & and_ln378_12_fu_9735_p2);

assign and_ln891_13_fu_10104_p2 = (tmp_157_fu_10052_p3 & and_ln378_13_fu_10046_p2);

assign and_ln891_14_fu_2662_p2 = (tmp_167_fu_2612_p3 & and_ln378_14_fu_2606_p2);

assign and_ln891_15_fu_4038_p2 = (tmp_173_reg_22579 & and_ln378_15_fu_4034_p2);

assign and_ln891_16_fu_4205_p2 = (tmp_179_fu_4153_p3 & and_ln378_16_fu_4147_p2);

assign and_ln891_17_fu_5064_p2 = (tmp_185_fu_5012_p3 & and_ln378_17_fu_5006_p2);

assign and_ln891_18_fu_6195_p2 = (tmp_195_reg_22808 & and_ln378_18_fu_6191_p2);

assign and_ln891_19_fu_6366_p2 = (tmp_201_fu_6314_p3 & and_ln378_19_fu_6308_p2);

assign and_ln891_1_fu_2454_p2 = (tmp_81_fu_2402_p3 & and_ln378_1_fu_2396_p2);

assign and_ln891_20_fu_7033_p2 = (tmp_207_fu_6981_p3 & and_ln378_20_fu_6975_p2);

assign and_ln891_21_fu_7767_p2 = (tmp_213_fu_7715_p3 & and_ln378_21_fu_7709_p2);

assign and_ln891_22_fu_8556_p2 = (tmp_221_fu_8504_p3 & and_ln378_22_fu_8498_p2);

assign and_ln891_23_fu_9236_p2 = (tmp_231_fu_9184_p3 & and_ln378_23_fu_9178_p2);

assign and_ln891_24_fu_2855_p2 = (tmp_239_fu_2805_p3 & and_ln378_24_fu_2799_p2);

assign and_ln891_25_fu_4273_p2 = (tmp_245_reg_22615 & and_ln378_25_fu_4269_p2);

assign and_ln891_26_fu_6437_p2 = (tmp_259_reg_22860 & and_ln378_26_fu_6433_p2);

assign and_ln891_27_fu_6608_p2 = (tmp_265_fu_6556_p3 & and_ln378_27_fu_6550_p2);

assign and_ln891_28_fu_7838_p2 = (tmp_275_reg_22987 & and_ln378_28_fu_7834_p2);

assign and_ln891_29_fu_8620_p2 = (tmp_285_reg_23053 & and_ln378_29_fu_8616_p2);

assign and_ln891_2_fu_3203_p2 = (tmp_87_fu_3151_p3 & and_ln378_2_fu_3145_p2);

assign and_ln891_30_fu_10480_p2 = (tmp_297_fu_10430_p3 & and_ln378_30_fu_10424_p2);

assign and_ln891_31_fu_11043_p2 = (tmp_303_fu_10991_p3 & and_ln378_31_fu_10985_p2);

assign and_ln891_32_fu_11718_p2 = (tmp_309_fu_11666_p3 & and_ln378_32_fu_11660_p2);

assign and_ln891_33_fu_10670_p2 = (tmp_315_fu_10620_p3 & and_ln378_33_fu_10614_p2);

assign and_ln891_34_fu_11273_p2 = (tmp_321_fu_11221_p3 & and_ln378_34_fu_11215_p2);

assign and_ln891_35_fu_11914_p2 = (tmp_327_fu_11862_p3 & and_ln378_35_fu_11856_p2);

assign and_ln891_36_fu_10844_p2 = (tmp_333_fu_10794_p3 & and_ln378_36_fu_10788_p2);

assign and_ln891_37_fu_11522_p2 = (tmp_339_fu_11470_p3 & and_ln378_37_fu_11464_p2);

assign and_ln891_38_fu_12120_p2 = (tmp_345_fu_12068_p3 & and_ln378_38_fu_12062_p2);

assign and_ln891_39_fu_13221_p2 = (tmp_351_fu_13171_p3 & and_ln378_39_fu_13165_p2);

assign and_ln891_3_fu_3956_p2 = (tmp_93_fu_3904_p3 & and_ln378_3_fu_3898_p2);

assign and_ln891_40_fu_13395_p2 = (tmp_361_fu_13345_p3 & and_ln378_40_fu_13339_p2);

assign and_ln891_41_fu_13565_p2 = (tmp_371_fu_13515_p3 & and_ln378_41_fu_13509_p2);

assign and_ln891_42_fu_17139_p2 = (tmp_377_reg_23624 & and_ln378_42_fu_17135_p2);

assign and_ln891_43_fu_13755_p2 = (tmp_385_fu_13705_p3 & and_ln378_43_fu_13699_p2);

assign and_ln891_44_fu_17227_p2 = (tmp_391_reg_23660 & and_ln378_44_fu_17223_p2);

assign and_ln891_45_fu_13929_p2 = (tmp_399_fu_13879_p3 & and_ln378_45_fu_13873_p2);

assign and_ln891_46_fu_15657_p2 = (tmp_405_fu_15605_p3 & and_ln378_46_fu_15599_p2);

assign and_ln891_47_fu_17443_p2 = (tmp_411_fu_17391_p3 & and_ln378_47_fu_17385_p2);

assign and_ln891_48_fu_14126_p2 = (tmp_417_fu_14076_p3 & and_ln378_48_fu_14070_p2);

assign and_ln891_49_fu_15894_p2 = (tmp_423_fu_15842_p3 & and_ln378_49_fu_15836_p2);

assign and_ln891_4_fu_4797_p2 = (tmp_99_fu_4745_p3 & and_ln378_4_fu_4739_p2);

assign and_ln891_50_fu_17655_p2 = (tmp_429_fu_17603_p3 & and_ln378_50_fu_17597_p2);

assign and_ln891_51_fu_16087_p2 = (tmp_435_fu_16037_p3 & and_ln378_51_fu_16031_p2);

assign and_ln891_52_fu_16261_p2 = (tmp_445_fu_16211_p3 & and_ln378_52_fu_16205_p2);

assign and_ln891_53_fu_14303_p2 = (tmp_455_fu_14253_p3 & and_ln378_53_fu_14247_p2);

assign and_ln891_54_fu_17967_p2 = (tmp_461_reg_23758 & and_ln378_54_fu_17963_p2);

assign and_ln891_55_fu_14493_p2 = (tmp_469_fu_14443_p3 & and_ln378_55_fu_14437_p2);

assign and_ln891_56_fu_18055_p2 = (tmp_475_reg_23794 & and_ln378_56_fu_18051_p2);

assign and_ln891_57_fu_14667_p2 = (tmp_483_fu_14617_p3 & and_ln378_57_fu_14611_p2);

assign and_ln891_58_fu_16815_p2 = (tmp_489_fu_16763_p3 & and_ln378_58_fu_16757_p2);

assign and_ln891_59_fu_18271_p2 = (tmp_495_fu_18219_p3 & and_ln378_59_fu_18213_p2);

assign and_ln891_5_fu_5418_p2 = (tmp_105_fu_5366_p3 & and_ln378_5_fu_5360_p2);

assign and_ln891_60_fu_14864_p2 = (tmp_501_fu_14814_p3 & and_ln378_60_fu_14808_p2);

assign and_ln891_61_fu_17052_p2 = (tmp_507_fu_17000_p3 & and_ln378_61_fu_16994_p2);

assign and_ln891_62_fu_18483_p2 = (tmp_513_fu_18431_p3 & and_ln378_62_fu_18425_p2);

assign and_ln891_6_fu_6108_p2 = (tmp_111_fu_6056_p3 & and_ln378_6_fu_6050_p2);

assign and_ln891_7_fu_6804_p2 = (tmp_117_fu_6752_p3 & and_ln378_7_fu_6746_p2);

assign and_ln891_8_fu_7516_p2 = (tmp_123_fu_7464_p3 & and_ln378_8_fu_7458_p2);

assign and_ln891_9_fu_8309_p2 = (tmp_129_fu_8257_p3 & and_ln378_9_fu_8251_p2);

assign and_ln891_fu_2087_p2 = (tmp_75_fu_2037_p3 & and_ln378_fu_2031_p2);

assign and_ln895_100_fu_15134_p2 = (xor_ln895_133_fu_15128_p2 & tmp_366_fu_15120_p3);

assign and_ln895_101_fu_13589_p2 = (xor_ln895_135_fu_13583_p2 & or_ln895_41_fu_13577_p2);

assign and_ln895_102_fu_15315_p2 = (xor_ln895_137_fu_15309_p2 & or_ln895_42_fu_15303_p2);

assign and_ln895_103_fu_17195_p2 = (xor_ln895_138_fu_17189_p2 & tmp_380_fu_17181_p3);

assign and_ln895_104_fu_13779_p2 = (xor_ln895_140_fu_13773_p2 & or_ln895_43_fu_13767_p2);

assign and_ln895_105_fu_15507_p2 = (xor_ln895_142_fu_15501_p2 & or_ln895_44_fu_15495_p2);

assign and_ln895_106_fu_17283_p2 = (xor_ln895_143_fu_17277_p2 & tmp_394_fu_17269_p3);

assign and_ln895_107_fu_13953_p2 = (xor_ln895_145_fu_13947_p2 & or_ln895_45_fu_13941_p2);

assign and_ln895_108_fu_15681_p2 = (xor_ln895_147_fu_15675_p2 & or_ln895_46_fu_15669_p2);

assign and_ln895_109_fu_17467_p2 = (xor_ln895_149_fu_17461_p2 & or_ln895_47_fu_17455_p2);

assign and_ln895_110_fu_14150_p2 = (xor_ln895_151_fu_14144_p2 & or_ln895_48_fu_14138_p2);

assign and_ln895_111_fu_15918_p2 = (xor_ln895_153_fu_15912_p2 & or_ln895_49_fu_15906_p2);

assign and_ln895_112_fu_17679_p2 = (xor_ln895_155_fu_17673_p2 & or_ln895_50_fu_17667_p2);

assign and_ln895_113_fu_16111_p2 = (xor_ln895_157_fu_16105_p2 & or_ln895_51_fu_16099_p2);

assign and_ln895_114_fu_17766_p2 = (xor_ln895_158_fu_17760_p2 & tmp_438_fu_17752_p3);

assign and_ln895_115_fu_17816_p2 = (xor_ln895_159_fu_17810_p2 & tmp_440_fu_17802_p3);

assign and_ln895_116_fu_16285_p2 = (xor_ln895_161_fu_16279_p2 & or_ln895_52_fu_16273_p2);

assign and_ln895_117_fu_17884_p2 = (xor_ln895_162_fu_17878_p2 & tmp_448_fu_17870_p3);

assign and_ln895_118_fu_17934_p2 = (xor_ln895_163_fu_17928_p2 & tmp_450_fu_17920_p3);

assign and_ln895_119_fu_14327_p2 = (xor_ln895_165_fu_14321_p2 & or_ln895_53_fu_14315_p2);

assign and_ln895_120_fu_16473_p2 = (xor_ln895_167_fu_16467_p2 & or_ln895_54_fu_16461_p2);

assign and_ln895_121_fu_18023_p2 = (xor_ln895_168_fu_18017_p2 & tmp_464_fu_18009_p3);

assign and_ln895_122_fu_14517_p2 = (xor_ln895_170_fu_14511_p2 & or_ln895_55_fu_14505_p2);

assign and_ln895_123_fu_16665_p2 = (xor_ln895_172_fu_16659_p2 & or_ln895_56_fu_16653_p2);

assign and_ln895_124_fu_18111_p2 = (xor_ln895_173_fu_18105_p2 & tmp_478_fu_18097_p3);

assign and_ln895_125_fu_14691_p2 = (xor_ln895_175_fu_14685_p2 & or_ln895_57_fu_14679_p2);

assign and_ln895_126_fu_16839_p2 = (xor_ln895_177_fu_16833_p2 & or_ln895_58_fu_16827_p2);

assign and_ln895_127_fu_18295_p2 = (xor_ln895_179_fu_18289_p2 & or_ln895_59_fu_18283_p2);

assign and_ln895_128_fu_14888_p2 = (xor_ln895_181_fu_14882_p2 & or_ln895_60_fu_14876_p2);

assign and_ln895_129_fu_17076_p2 = (xor_ln895_183_fu_17070_p2 & or_ln895_61_fu_17064_p2);

assign and_ln895_130_fu_18507_p2 = (xor_ln895_185_fu_18501_p2 & or_ln895_62_fu_18495_p2);

assign and_ln895_131_fu_12262_p2 = (xor_ln895_186_fu_12256_p2 & tmp_516_fu_12248_p3);

assign and_ln895_132_fu_12312_p2 = (xor_ln895_187_fu_12306_p2 & tmp_518_fu_12298_p3);

assign and_ln895_133_fu_12362_p2 = (xor_ln895_188_fu_12356_p2 & tmp_520_fu_12348_p3);

assign and_ln895_134_fu_12427_p2 = (xor_ln895_189_fu_12421_p2 & or_ln895_63_fu_12415_p2);

assign and_ln895_135_fu_12495_p2 = (xor_ln895_190_fu_12489_p2 & tmp_525_fu_12481_p3);

assign and_ln895_136_fu_12584_p2 = (xor_ln895_191_fu_12578_p2 & or_ln895_64_fu_12572_p2);

assign and_ln895_137_fu_12694_p2 = (xor_ln895_192_fu_12688_p2 & or_ln895_65_fu_12682_p2);

assign and_ln895_138_fu_12762_p2 = (xor_ln895_193_fu_12756_p2 & tmp_533_fu_12748_p3);

assign and_ln895_139_fu_12812_p2 = (xor_ln895_194_fu_12806_p2 & tmp_535_fu_12798_p3);

assign and_ln895_140_fu_12915_p2 = (xor_ln895_195_fu_12909_p2 & or_ln895_66_fu_12903_p2);

assign and_ln895_141_fu_12983_p2 = (xor_ln895_196_fu_12977_p2 & tmp_540_fu_12969_p3);

assign and_ln895_142_fu_13064_p2 = (xor_ln895_197_fu_13058_p2 & or_ln895_67_fu_13052_p2);

assign and_ln895_143_fu_18601_p2 = (xor_ln895_198_fu_18595_p2 & tmp_545_fu_18587_p3);

assign and_ln895_144_fu_18672_p2 = (xor_ln895_199_fu_18666_p2 & tmp_547_fu_18658_p3);

assign and_ln895_145_fu_18777_p2 = (xor_ln895_200_fu_18771_p2 & tmp_549_fu_18763_p3);

assign and_ln895_146_fu_18848_p2 = (xor_ln895_201_fu_18842_p2 & tmp_551_fu_18834_p3);

assign and_ln895_147_fu_18953_p2 = (xor_ln895_202_fu_18947_p2 & tmp_553_fu_18939_p3);

assign and_ln895_148_fu_19024_p2 = (xor_ln895_203_fu_19018_p2 & tmp_555_fu_19010_p3);

assign and_ln895_149_fu_19129_p2 = (xor_ln895_204_fu_19123_p2 & tmp_557_fu_19115_p3);

assign and_ln895_150_fu_19200_p2 = (xor_ln895_205_fu_19194_p2 & tmp_559_fu_19186_p3);

assign and_ln895_151_fu_19305_p2 = (xor_ln895_206_fu_19299_p2 & tmp_561_fu_19291_p3);

assign and_ln895_152_fu_19376_p2 = (xor_ln895_207_fu_19370_p2 & tmp_563_fu_19362_p3);

assign and_ln895_153_fu_19481_p2 = (xor_ln895_208_fu_19475_p2 & tmp_565_fu_19467_p3);

assign and_ln895_154_fu_19552_p2 = (xor_ln895_209_fu_19546_p2 & tmp_567_fu_19538_p3);

assign and_ln895_155_fu_19657_p2 = (xor_ln895_210_fu_19651_p2 & tmp_569_fu_19643_p3);

assign and_ln895_156_fu_19728_p2 = (xor_ln895_211_fu_19722_p2 & tmp_571_fu_19714_p3);

assign and_ln895_157_fu_19833_p2 = (xor_ln895_212_fu_19827_p2 & tmp_573_fu_19819_p3);

assign and_ln895_158_fu_19904_p2 = (xor_ln895_213_fu_19898_p2 & tmp_575_fu_19890_p3);

assign and_ln895_159_fu_20009_p2 = (xor_ln895_214_fu_20003_p2 & tmp_577_fu_19995_p3);

assign and_ln895_160_fu_20080_p2 = (xor_ln895_215_fu_20074_p2 & tmp_579_fu_20066_p3);

assign and_ln895_161_fu_20183_p2 = (xor_ln895_216_fu_20177_p2 & tmp_581_fu_20169_p3);

assign and_ln895_162_fu_20252_p2 = (xor_ln895_217_fu_20246_p2 & tmp_583_fu_20238_p3);

assign and_ln895_163_fu_20321_p2 = (xor_ln895_218_fu_20315_p2 & tmp_585_fu_20307_p3);

assign and_ln895_164_fu_20390_p2 = (xor_ln895_219_fu_20384_p2 & tmp_587_fu_20376_p3);

assign and_ln895_165_fu_20459_p2 = (xor_ln895_220_fu_20453_p2 & tmp_589_fu_20445_p3);

assign and_ln895_166_fu_20528_p2 = (xor_ln895_221_fu_20522_p2 & tmp_591_fu_20514_p3);

assign and_ln895_167_fu_20597_p2 = (xor_ln895_222_fu_20591_p2 & tmp_593_fu_20583_p3);

assign and_ln895_168_fu_20666_p2 = (xor_ln895_223_fu_20660_p2 & tmp_595_fu_20652_p3);

assign and_ln895_169_fu_20735_p2 = (xor_ln895_224_fu_20729_p2 & tmp_597_fu_20721_p3);

assign and_ln895_170_fu_20804_p2 = (xor_ln895_225_fu_20798_p2 & tmp_599_fu_20790_p3);

assign and_ln895_171_fu_20873_p2 = (xor_ln895_226_fu_20867_p2 & tmp_601_fu_20859_p3);

assign and_ln895_172_fu_20942_p2 = (xor_ln895_227_fu_20936_p2 & tmp_603_fu_20928_p3);

assign and_ln895_173_fu_21011_p2 = (xor_ln895_228_fu_21005_p2 & tmp_605_fu_20997_p3);

assign and_ln895_174_fu_21080_p2 = (xor_ln895_229_fu_21074_p2 & tmp_607_fu_21066_p3);

assign and_ln895_175_fu_21149_p2 = (xor_ln895_230_fu_21143_p2 & tmp_609_fu_21135_p3);

assign and_ln895_176_fu_21218_p2 = (xor_ln895_231_fu_21212_p2 & tmp_611_fu_21204_p3);

assign and_ln895_177_fu_21287_p2 = (xor_ln895_232_fu_21281_p2 & tmp_613_fu_21273_p3);

assign and_ln895_178_fu_21356_p2 = (xor_ln895_233_fu_21350_p2 & tmp_615_fu_21342_p3);

assign and_ln895_18_fu_1421_p2 = (xor_ln895_18_fu_1415_p2 & tmp_38_fu_1407_p3);

assign and_ln895_19_fu_1499_p2 = (xor_ln895_19_fu_1493_p2 & tmp_40_fu_1485_p3);

assign and_ln895_20_fu_1651_p2 = (xor_ln895_20_fu_1645_p2 & tmp_42_fu_1637_p3);

assign and_ln895_21_fu_1569_p2 = (xor_ln895_21_fu_1563_p2 & tmp_44_fu_1555_p3);

assign and_ln895_22_fu_1721_p2 = (xor_ln895_22_fu_1715_p2 & tmp_46_fu_1707_p3);

assign and_ln895_23_fu_1879_p2 = (xor_ln895_23_fu_1873_p2 & tmp_48_fu_1865_p3);

assign and_ln895_24_fu_1949_p2 = (xor_ln895_24_fu_1943_p2 & tmp_50_fu_1935_p3);

assign and_ln895_25_fu_2220_p2 = (xor_ln895_25_fu_2214_p2 & tmp_52_fu_2206_p3);

assign and_ln895_26_fu_2290_p2 = (xor_ln895_26_fu_2284_p2 & tmp_54_fu_2276_p3);

assign and_ln895_27_fu_2973_p2 = (xor_ln895_10_fu_2967_p2 & tmp_56_fu_2959_p3);

assign and_ln895_28_fu_3043_p2 = (xor_ln895_11_fu_3037_p2 & tmp_58_fu_3029_p3);

assign and_ln895_29_fu_3692_p2 = (xor_ln895_12_fu_3686_p2 & tmp_60_fu_3678_p3);

assign and_ln895_30_fu_3762_p2 = (xor_ln895_13_fu_3756_p2 & tmp_62_fu_3748_p3);

assign and_ln895_31_fu_4549_p2 = (xor_ln895_14_fu_4543_p2 & tmp_64_fu_4535_p3);

assign and_ln895_32_fu_4619_p2 = (xor_ln895_15_fu_4613_p2 & tmp_66_fu_4605_p3);

assign and_ln895_33_fu_5184_p2 = (xor_ln895_16_fu_5178_p2 & tmp_68_fu_5170_p3);

assign and_ln895_34_fu_5254_p2 = (xor_ln895_17_fu_5248_p2 & tmp_70_fu_5240_p3);

assign and_ln895_35_fu_2111_p2 = (xor_ln895_28_fu_2105_p2 & or_ln895_fu_2099_p2);

assign and_ln895_36_fu_2478_p2 = (xor_ln895_30_fu_2472_p2 & or_ln895_1_fu_2466_p2);

assign and_ln895_37_fu_3227_p2 = (xor_ln895_32_fu_3221_p2 & or_ln895_2_fu_3215_p2);

assign and_ln895_38_fu_3980_p2 = (xor_ln895_34_fu_3974_p2 & or_ln895_3_fu_3968_p2);

assign and_ln895_39_fu_4821_p2 = (xor_ln895_36_fu_4815_p2 & or_ln895_4_fu_4809_p2);

assign and_ln895_40_fu_5442_p2 = (xor_ln895_38_fu_5436_p2 & or_ln895_5_fu_5430_p2);

assign and_ln895_41_fu_6132_p2 = (xor_ln895_40_fu_6126_p2 & or_ln895_6_fu_6120_p2);

assign and_ln895_42_fu_6828_p2 = (xor_ln895_42_fu_6822_p2 & or_ln895_7_fu_6816_p2);

assign and_ln895_43_fu_7540_p2 = (xor_ln895_44_fu_7534_p2 & or_ln895_8_fu_7528_p2);

assign and_ln895_44_fu_8333_p2 = (xor_ln895_46_fu_8327_p2 & or_ln895_9_fu_8321_p2);

assign and_ln895_45_fu_8947_p2 = (xor_ln895_48_fu_8941_p2 & or_ln895_10_fu_8935_p2);

assign and_ln895_46_fu_9456_p2 = (xor_ln895_50_fu_9450_p2 & or_ln895_11_fu_9444_p2);

assign and_ln895_47_fu_9817_p2 = (xor_ln895_52_fu_9811_p2 & or_ln895_12_fu_9805_p2);

assign and_ln895_48_fu_9902_p2 = (xor_ln895_53_fu_9896_p2 & tmp_150_fu_9888_p3);

assign and_ln895_49_fu_9952_p2 = (xor_ln895_54_fu_9946_p2 & tmp_152_fu_9938_p3);

assign and_ln895_50_fu_10128_p2 = (xor_ln895_56_fu_10122_p2 & or_ln895_13_fu_10116_p2);

assign and_ln895_51_fu_10199_p2 = (xor_ln895_57_fu_10193_p2 & tmp_160_fu_10185_p3);

assign and_ln895_52_fu_10249_p2 = (xor_ln895_58_fu_10243_p2 & tmp_162_fu_10235_p3);

assign and_ln895_53_fu_2686_p2 = (xor_ln895_60_fu_2680_p2 & or_ln895_14_fu_2674_p2);

assign and_ln895_54_fu_3458_p2 = (xor_ln895_62_fu_3452_p2 & or_ln895_15_fu_3446_p2);

assign and_ln895_55_fu_4229_p2 = (xor_ln895_64_fu_4223_p2 & or_ln895_16_fu_4217_p2);

assign and_ln895_56_fu_5088_p2 = (xor_ln895_66_fu_5082_p2 & or_ln895_17_fu_5076_p2);

assign and_ln895_57_fu_5543_p2 = (xor_ln895_67_fu_5537_p2 & tmp_188_fu_5529_p3);

assign and_ln895_58_fu_5593_p2 = (xor_ln895_68_fu_5587_p2 & tmp_190_fu_5579_p3);

assign and_ln895_59_fu_5766_p2 = (xor_ln895_70_fu_5760_p2 & or_ln895_18_fu_5754_p2);

assign and_ln895_60_fu_6390_p2 = (xor_ln895_72_fu_6384_p2 & or_ln895_19_fu_6378_p2);

assign and_ln895_61_fu_7057_p2 = (xor_ln895_74_fu_7051_p2 & or_ln895_20_fu_7045_p2);

assign and_ln895_62_fu_7791_p2 = (xor_ln895_76_fu_7785_p2 & or_ln895_21_fu_7779_p2);

assign and_ln895_63_fu_8404_p2 = (xor_ln895_77_fu_8398_p2 & tmp_216_fu_8390_p3);

assign and_ln895_64_fu_8580_p2 = (xor_ln895_79_fu_8574_p2 & or_ln895_22_fu_8568_p2);

assign and_ln895_65_fu_9034_p2 = (xor_ln895_80_fu_9028_p2 & tmp_224_fu_9020_p3);

assign and_ln895_66_fu_9084_p2 = (xor_ln895_81_fu_9078_p2 & tmp_226_fu_9070_p3);

assign and_ln895_67_fu_9260_p2 = (xor_ln895_83_fu_9254_p2 & or_ln895_23_fu_9248_p2);

assign and_ln895_68_fu_9527_p2 = (xor_ln895_84_fu_9521_p2 & tmp_234_fu_9513_p3);

assign and_ln895_69_fu_2879_p2 = (xor_ln895_86_fu_2873_p2 & or_ln895_24_fu_2867_p2);

assign and_ln895_70_fu_3632_p2 = (xor_ln895_88_fu_3626_p2 & or_ln895_25_fu_3620_p2);

assign and_ln895_71_fu_4329_p2 = (xor_ln895_89_fu_4323_p2 & tmp_248_fu_4315_p3);

assign and_ln895_72_fu_4379_p2 = (xor_ln895_90_fu_4373_p2 & tmp_250_fu_4365_p3);

assign and_ln895_73_fu_4429_p2 = (xor_ln895_91_fu_4423_p2 & tmp_252_fu_4415_p3);

assign and_ln895_74_fu_4479_p2 = (xor_ln895_92_fu_4473_p2 & tmp_254_fu_4465_p3);

assign and_ln895_75_fu_5947_p2 = (xor_ln895_94_fu_5941_p2 & or_ln895_26_fu_5935_p2);

assign and_ln895_76_fu_6632_p2 = (xor_ln895_96_fu_6626_p2 & or_ln895_27_fu_6620_p2);

assign and_ln895_77_fu_7144_p2 = (xor_ln895_97_fu_7138_p2 & tmp_268_fu_7130_p3);

assign and_ln895_78_fu_7194_p2 = (xor_ln895_98_fu_7188_p2 & tmp_270_fu_7180_p3);

assign and_ln895_79_fu_7366_p2 = (xor_ln895_100_fu_7360_p2 & or_ln895_28_fu_7354_p2);

assign and_ln895_80_fu_7894_p2 = (xor_ln895_101_fu_7888_p2 & tmp_278_fu_7880_p3);

assign and_ln895_81_fu_7944_p2 = (xor_ln895_102_fu_7938_p2 & tmp_280_fu_7930_p3);

assign and_ln895_82_fu_8116_p2 = (xor_ln895_104_fu_8110_p2 & or_ln895_29_fu_8104_p2);

assign and_ln895_83_fu_10312_p2 = (xor_ln895_105_fu_10306_p2 & tmp_288_fu_10298_p3);

assign and_ln895_84_fu_9590_p2 = (xor_ln895_106_fu_9584_p2 & tmp_290_fu_9576_p3);

assign and_ln895_85_fu_8689_p2 = (xor_ln895_107_fu_8683_p2 & tmp_292_fu_8675_p3);

assign and_ln895_86_fu_10504_p2 = (xor_ln895_109_fu_10498_p2 & or_ln895_30_fu_10492_p2);

assign and_ln895_87_fu_11067_p2 = (xor_ln895_111_fu_11061_p2 & or_ln895_31_fu_11055_p2);

assign and_ln895_88_fu_11742_p2 = (xor_ln895_113_fu_11736_p2 & or_ln895_32_fu_11730_p2);

assign and_ln895_89_fu_10694_p2 = (xor_ln895_115_fu_10688_p2 & or_ln895_33_fu_10682_p2);

assign and_ln895_90_fu_11297_p2 = (xor_ln895_117_fu_11291_p2 & or_ln895_34_fu_11285_p2);

assign and_ln895_91_fu_11938_p2 = (xor_ln895_119_fu_11932_p2 & or_ln895_35_fu_11926_p2);

assign and_ln895_92_fu_10868_p2 = (xor_ln895_121_fu_10862_p2 & or_ln895_36_fu_10856_p2);

assign and_ln895_93_fu_11546_p2 = (xor_ln895_123_fu_11540_p2 & or_ln895_37_fu_11534_p2);

assign and_ln895_94_fu_12144_p2 = (xor_ln895_125_fu_12138_p2 & or_ln895_38_fu_12132_p2);

assign and_ln895_95_fu_13245_p2 = (xor_ln895_127_fu_13239_p2 & or_ln895_39_fu_13233_p2);

assign and_ln895_96_fu_14966_p2 = (xor_ln895_128_fu_14960_p2 & tmp_354_fu_14952_p3);

assign and_ln895_97_fu_15016_p2 = (xor_ln895_129_fu_15010_p2 & tmp_356_fu_15002_p3);

assign and_ln895_98_fu_13419_p2 = (xor_ln895_131_fu_13413_p2 & or_ln895_40_fu_13407_p2);

assign and_ln895_99_fu_15084_p2 = (xor_ln895_132_fu_15078_p2 & tmp_364_fu_15070_p3);

assign and_ln895_fu_1351_p2 = (xor_ln895_fu_1345_p2 & tmp_36_fu_1337_p3);

assign and_ln896_10_fu_8971_p2 = (xor_ln896_62_fu_8965_p2 & tmp_131_fu_8816_p3);

assign and_ln896_11_fu_9480_p2 = (xor_ln896_63_fu_9474_p2 & tmp_137_fu_9325_p3);

assign and_ln896_12_fu_9841_p2 = (xor_ln896_64_fu_9835_p2 & tmp_143_fu_9686_p3);

assign and_ln896_13_fu_10152_p2 = (xor_ln896_65_fu_10146_p2 & tmp_153_fu_9997_p3);

assign and_ln896_14_fu_2710_p2 = (xor_ln896_70_fu_2704_p2 & tmp_163_fu_2552_p3);

assign and_ln896_15_fu_4048_p2 = (xor_ln896_71_fu_4043_p2 & tmp_169_reg_22559);

assign and_ln896_16_fu_4253_p2 = (xor_ln896_74_fu_4247_p2 & tmp_175_fu_4098_p3);

assign and_ln896_17_fu_5112_p2 = (xor_ln896_75_fu_5106_p2 & tmp_181_fu_4957_p3);

assign and_ln896_18_fu_6205_p2 = (xor_ln896_98_fu_6200_p2 & tmp_191_reg_22788);

assign and_ln896_19_fu_6414_p2 = (xor_ln896_99_fu_6408_p2 & tmp_197_fu_6259_p3);

assign and_ln896_1_fu_2502_p2 = (xor_ln896_27_fu_2496_p2 & tmp_77_fu_2347_p3);

assign and_ln896_20_fu_7081_p2 = (xor_ln896_102_fu_7075_p2 & tmp_203_fu_6926_p3);

assign and_ln896_21_fu_7815_p2 = (xor_ln896_103_fu_7809_p2 & tmp_209_fu_7651_p3);

assign and_ln896_22_fu_8604_p2 = (xor_ln896_108_fu_8598_p2 & tmp_217_fu_8449_p3);

assign and_ln896_23_fu_9284_p2 = (xor_ln896_113_fu_9278_p2 & tmp_227_fu_9129_p3);

assign and_ln896_24_fu_2903_p2 = (xor_ln896_128_fu_2897_p2 & tmp_235_fu_2745_p3);

assign and_ln896_25_fu_4283_p2 = (xor_ln896_129_fu_4278_p2 & tmp_241_reg_22595);

assign and_ln896_26_fu_6447_p2 = (xor_ln896_132_fu_6442_p2 & tmp_255_reg_22840);

assign and_ln896_27_fu_6656_p2 = (xor_ln896_133_fu_6650_p2 & tmp_261_fu_6501_p3);

assign and_ln896_28_fu_7848_p2 = (xor_ln896_138_fu_7843_p2 & tmp_271_reg_22967);

assign and_ln896_29_fu_8630_p2 = (xor_ln896_143_fu_8625_p2 & tmp_281_reg_23033);

assign and_ln896_2_fu_3251_p2 = (xor_ln896_30_fu_3245_p2 & tmp_83_fu_3096_p3);

assign and_ln896_30_fu_10528_p2 = (xor_ln896_156_fu_10522_p2 & tmp_293_fu_10366_p3);

assign and_ln896_31_fu_11091_p2 = (xor_ln896_157_fu_11085_p2 & tmp_299_fu_10936_p3);

assign and_ln896_32_fu_11766_p2 = (xor_ln896_158_fu_11760_p2 & tmp_305_fu_11611_p3);

assign and_ln896_33_fu_10718_p2 = (xor_ln896_160_fu_10712_p2 & tmp_311_fu_10556_p3);

assign and_ln896_34_fu_11321_p2 = (xor_ln896_162_fu_11315_p2 & tmp_317_fu_11166_p3);

assign and_ln896_35_fu_11962_p2 = (xor_ln896_163_fu_11956_p2 & tmp_323_fu_11807_p3);

assign and_ln896_36_fu_10892_p2 = (xor_ln896_164_fu_10886_p2 & tmp_329_fu_10730_p3);

assign and_ln896_37_fu_11570_p2 = (xor_ln896_165_fu_11564_p2 & tmp_335_fu_11415_p3);

assign and_ln896_38_fu_12168_p2 = (xor_ln896_166_fu_12162_p2 & tmp_341_fu_12013_p3);

assign and_ln896_39_fu_13269_p2 = (xor_ln896_167_fu_13263_p2 & tmp_347_fu_13111_p3);

assign and_ln896_3_fu_4004_p2 = (xor_ln896_31_fu_3998_p2 & tmp_89_fu_3849_p3);

assign and_ln896_40_fu_13443_p2 = (xor_ln896_168_fu_13437_p2 & tmp_357_fu_13281_p3);

assign and_ln896_41_fu_13613_p2 = (xor_ln896_169_fu_13607_p2 & tmp_367_fu_13455_p3);

assign and_ln896_42_fu_17149_p2 = (xor_ln896_170_fu_17144_p2 & tmp_373_reg_23604);

assign and_ln896_43_fu_13803_p2 = (xor_ln896_171_fu_13797_p2 & tmp_381_fu_13641_p3);

assign and_ln896_44_fu_17237_p2 = (xor_ln896_172_fu_17232_p2 & tmp_387_reg_23640);

assign and_ln896_45_fu_13977_p2 = (xor_ln896_173_fu_13971_p2 & tmp_395_fu_13815_p3);

assign and_ln896_46_fu_15705_p2 = (xor_ln896_174_fu_15699_p2 & tmp_401_fu_15550_p3);

assign and_ln896_47_fu_17491_p2 = (xor_ln896_175_fu_17485_p2 & tmp_407_fu_17336_p3);

assign and_ln896_48_fu_14174_p2 = (xor_ln896_176_fu_14168_p2 & tmp_413_fu_14012_p3);

assign and_ln896_49_fu_15942_p2 = (xor_ln896_177_fu_15936_p2 & tmp_419_fu_15787_p3);

assign and_ln896_4_fu_4845_p2 = (xor_ln896_40_fu_4839_p2 & tmp_95_fu_4690_p3);

assign and_ln896_50_fu_17703_p2 = (xor_ln896_178_fu_17697_p2 & tmp_425_fu_17548_p3);

assign and_ln896_51_fu_16135_p2 = (xor_ln896_179_fu_16129_p2 & tmp_431_fu_15977_p3);

assign and_ln896_52_fu_16309_p2 = (xor_ln896_180_fu_16303_p2 & tmp_441_fu_16147_p3);

assign and_ln896_53_fu_14351_p2 = (xor_ln896_181_fu_14345_p2 & tmp_451_fu_14193_p3);

assign and_ln896_54_fu_17977_p2 = (xor_ln896_182_fu_17972_p2 & tmp_457_reg_23738);

assign and_ln896_55_fu_14541_p2 = (xor_ln896_183_fu_14535_p2 & tmp_465_fu_14379_p3);

assign and_ln896_56_fu_18065_p2 = (xor_ln896_184_fu_18060_p2 & tmp_471_reg_23774);

assign and_ln896_57_fu_14715_p2 = (xor_ln896_185_fu_14709_p2 & tmp_479_fu_14553_p3);

assign and_ln896_58_fu_16863_p2 = (xor_ln896_186_fu_16857_p2 & tmp_485_fu_16708_p3);

assign and_ln896_59_fu_18319_p2 = (xor_ln896_187_fu_18313_p2 & tmp_491_fu_18164_p3);

assign and_ln896_5_fu_5466_p2 = (xor_ln896_41_fu_5460_p2 & tmp_101_fu_5311_p3);

assign and_ln896_60_fu_14912_p2 = (xor_ln896_188_fu_14906_p2 & tmp_497_fu_14750_p3);

assign and_ln896_61_fu_17100_p2 = (xor_ln896_189_fu_17094_p2 & tmp_503_fu_16945_p3);

assign and_ln896_62_fu_18531_p2 = (xor_ln896_190_fu_18525_p2 & tmp_509_fu_18376_p3);

assign and_ln896_63_fu_12433_p2 = (tmp_523_fu_12407_p3 & tmp_522_fu_12399_p3);

assign and_ln896_64_fu_12445_p2 = (xor_ln896_159_fu_12439_p2 & tmp_521_fu_12391_p3);

assign and_ln896_65_fu_12590_p2 = (tmp_528_fu_12564_p3 & tmp_527_fu_12556_p3);

assign and_ln896_66_fu_12602_p2 = (xor_ln896_161_fu_12596_p2 & tmp_526_fu_12548_p3);

assign and_ln896_67_fu_12700_p2 = (tmp_531_fu_12674_p3 & tmp_530_fu_12666_p3);

assign and_ln896_68_fu_12712_p2 = (xor_ln896_191_fu_12706_p2 & tmp_529_fu_12648_p3);

assign and_ln896_69_fu_12921_p2 = (tmp_538_fu_12895_p3 & tmp_537_fu_12887_p3);

assign and_ln896_6_fu_6156_p2 = (xor_ln896_50_fu_6150_p2 & tmp_107_fu_6001_p3);

assign and_ln896_70_fu_12933_p2 = (xor_ln896_192_fu_12927_p2 & tmp_536_fu_12869_p3);

assign and_ln896_71_fu_13070_p2 = (tmp_543_fu_13044_p3 & tmp_542_fu_13036_p3);

assign and_ln896_72_fu_13082_p2 = (xor_ln896_193_fu_13076_p2 & tmp_541_fu_13018_p3);

assign and_ln896_7_fu_6852_p2 = (xor_ln896_53_fu_6846_p2 & tmp_113_fu_6697_p3);

assign and_ln896_8_fu_7564_p2 = (xor_ln896_54_fu_7558_p2 & tmp_119_fu_7409_p3);

assign and_ln896_9_fu_8357_p2 = (xor_ln896_57_fu_8351_p2 & tmp_125_fu_8193_p3);

assign and_ln896_fu_2135_p2 = (xor_ln896_26_fu_2129_p2 & tmp_71_fu_1977_p3);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];

assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];

assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];

assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];

assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];

assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];

assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];

assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];

assign ap_CS_fsm_state34 = ap_CS_fsm[32'd33];

assign ap_CS_fsm_state35 = ap_CS_fsm[32'd34];

assign ap_CS_fsm_state36 = ap_CS_fsm[32'd35];

assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];

assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];

assign ap_CS_fsm_state39 = ap_CS_fsm[32'd38];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state40 = ap_CS_fsm[32'd39];

assign ap_CS_fsm_state41 = ap_CS_fsm[32'd40];

assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];

assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];

assign ap_CS_fsm_state44 = ap_CS_fsm[32'd43];

assign ap_CS_fsm_state45 = ap_CS_fsm[32'd44];

assign ap_CS_fsm_state46 = ap_CS_fsm[32'd45];

assign ap_CS_fsm_state47 = ap_CS_fsm[32'd46];

assign ap_CS_fsm_state48 = ap_CS_fsm[32'd47];

assign ap_CS_fsm_state49 = ap_CS_fsm[32'd48];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state50 = ap_CS_fsm[32'd49];

assign ap_CS_fsm_state51 = ap_CS_fsm[32'd50];

assign ap_CS_fsm_state52 = ap_CS_fsm[32'd51];

assign ap_CS_fsm_state53 = ap_CS_fsm[32'd52];

assign ap_CS_fsm_state54 = ap_CS_fsm[32'd53];

assign ap_CS_fsm_state55 = ap_CS_fsm[32'd54];

assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];

assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];

assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];

assign ap_CS_fsm_state59 = ap_CS_fsm[32'd58];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state60 = ap_CS_fsm[32'd59];

assign ap_CS_fsm_state61 = ap_CS_fsm[32'd60];

assign ap_CS_fsm_state62 = ap_CS_fsm[32'd61];

assign ap_CS_fsm_state63 = ap_CS_fsm[32'd62];

assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];

assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];

assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];

assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];

assign ap_CS_fsm_state68 = ap_CS_fsm[32'd67];

assign ap_CS_fsm_state69 = ap_CS_fsm[32'd68];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];

assign ap_CS_fsm_state71 = ap_CS_fsm[32'd70];

assign ap_CS_fsm_state72 = ap_CS_fsm[32'd71];

assign ap_CS_fsm_state73 = ap_CS_fsm[32'd72];

assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];

assign ap_CS_fsm_state75 = ap_CS_fsm[32'd74];

assign ap_CS_fsm_state76 = ap_CS_fsm[32'd75];

assign ap_CS_fsm_state77 = ap_CS_fsm[32'd76];

assign ap_CS_fsm_state78 = ap_CS_fsm[32'd77];

assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

assign ap_CS_fsm_state81 = ap_CS_fsm[32'd80];

assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];

assign ap_CS_fsm_state83 = ap_CS_fsm[32'd82];

assign ap_CS_fsm_state84 = ap_CS_fsm[32'd83];

assign ap_CS_fsm_state85 = ap_CS_fsm[32'd84];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

assign ap_NS_fsm_state12 = ap_NS_fsm[32'd11];

assign ap_NS_fsm_state2 = ap_NS_fsm[32'd1];

assign ap_NS_fsm_state46 = ap_NS_fsm[32'd45];

assign ap_NS_fsm_state66 = ap_NS_fsm[32'd65];

assign ap_block_state10_pp0_stage9_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage10_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage11_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage12_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage13_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage14_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage15_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage16_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage17_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage18_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0 = (ap_start_int == 1'b0);
end

assign ap_block_state20_pp0_stage19_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage20_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage21_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage22_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage23_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state25_pp0_stage24_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state26_pp0_stage25_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state27_pp0_stage26_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state28_pp0_stage27_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state29_pp0_stage28_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state30_pp0_stage29_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state31_pp0_stage30_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state32_pp0_stage31_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state33_pp0_stage32_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state34_pp0_stage33_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state35_pp0_stage34_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state36_pp0_stage35_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state37_pp0_stage36_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state38_pp0_stage37_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state39_pp0_stage38_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state40_pp0_stage39_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state41_pp0_stage40_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state42_pp0_stage41_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state43_pp0_stage42_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state44_pp0_stage43_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state45_pp0_stage44_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state46_pp0_stage45_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state47_pp0_stage46_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state48_pp0_stage47_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state49_pp0_stage48_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state50_pp0_stage49_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state51_pp0_stage50_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state52_pp0_stage51_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state53_pp0_stage52_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state54_pp0_stage53_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state55_pp0_stage54_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state56_pp0_stage55_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state57_pp0_stage56_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state58_pp0_stage57_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state59_pp0_stage58_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage4_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state60_pp0_stage59_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state61_pp0_stage60_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state62_pp0_stage61_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state63_pp0_stage62_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state64_pp0_stage63_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state65_pp0_stage64_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state66_pp0_stage65_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state67_pp0_stage66_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state68_pp0_stage67_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state69_pp0_stage68_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage5_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state70_pp0_stage69_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state71_pp0_stage70_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state72_pp0_stage71_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state73_pp0_stage72_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state74_pp0_stage73_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state75_pp0_stage74_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state76_pp0_stage75_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state77_pp0_stage76_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state78_pp0_stage77_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state79_pp0_stage78_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage6_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state80_pp0_stage79_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state81_pp0_stage80_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state82_pp0_stage81_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state83_pp0_stage82_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state84_pp0_stage83_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state85_pp0_stage84_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage7_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage8_iter0 = ~(1'b1 == 1'b1);

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

assign grp_fu_1188_p2 = (($signed(temp5_q1) > $signed(21'd0)) ? 1'b1 : 1'b0);

assign grp_fu_1194_p2 = (($signed(temp5_q0) > $signed(21'd0)) ? 1'b1 : 1'b0);

assign grp_fu_21385_p1 = 35'd34359732525;

assign grp_fu_21397_p1 = 28'd268435419;

assign grp_fu_21404_p0 = sext_ln1273_2_fu_1597_p1;

assign grp_fu_21404_p1 = 35'd34359734235;

assign grp_fu_21411_p1 = 34'd17179866261;

assign grp_fu_21418_p0 = sext_ln1273_2_fu_1597_p1;

assign grp_fu_21418_p1 = 35'd34359732525;

assign grp_fu_21430_p0 = sext_ln1273_6_fu_1601_p1;

assign grp_fu_21430_p1 = 35'd34359734235;

assign grp_fu_21437_p0 = sext_ln1273_6_fu_1601_p1;

assign grp_fu_21437_p1 = 35'd34359732525;

assign grp_fu_21449_p1 = 30'd1073741686;

assign grp_fu_21456_p1 = 28'd268435419;

assign grp_fu_21465_p1 = 28'd268435419;

assign grp_fu_21474_p1 = 35'd5843;

assign grp_fu_21481_p1 = 28'd37;

assign grp_fu_21488_p0 = sext_ln1273_12_fu_2544_p1;

assign grp_fu_21488_p1 = 35'd4133;

assign grp_fu_21495_p0 = sext_ln1273_12_fu_2544_p1;

assign grp_fu_21495_p1 = 35'd5843;

assign grp_fu_21502_p1 = 28'd37;

assign grp_fu_21509_p1 = 34'd2923;

assign grp_fu_21516_p1 = 30'd138;

assign grp_fu_21523_p0 = sext_ln1273_16_fu_3286_p1;

assign grp_fu_21523_p1 = 35'd4133;

assign grp_fu_21530_p0 = sext_ln1273_16_fu_3286_p1;

assign grp_fu_21530_p1 = 35'd5843;

assign grp_fu_21539_p1 = 28'd37;

assign grp_fu_21546_p1 = 36'd68719463936;

assign grp_fu_21553_p1 = 36'd68719463936;

assign grp_fu_21560_p1 = 36'd12800;

assign grp_fu_21567_p1 = 36'd68719463936;

assign grp_fu_21575_p1 = 36'd12800;

assign grp_fu_21582_p1 = 36'd12800;

assign grp_fu_21590_p0 = sext_ln1273_37_fu_8721_p1;

assign grp_fu_21590_p1 = 30'd1073741649;

assign grp_fu_21597_p1 = 35'd4204;

assign grp_fu_21604_p1 = 31'd2147483290;

assign grp_fu_21611_p1 = 34'd4061;

assign grp_fu_21618_p1 = 34'd3973;

assign grp_fu_21630_p1 = 31'd2147483290;

assign grp_fu_21642_p1 = 30'd1073741649;

assign grp_fu_21654_p0 = sext_ln1273_44_fu_12228_p1;

assign grp_fu_21654_p1 = 35'd7479;

assign grp_fu_21666_p1 = 28'd47;

assign grp_fu_21678_p0 = sext_ln1273_44_fu_12228_p1;

assign grp_fu_21678_p1 = 35'd5290;

assign grp_fu_21690_p0 = sext_ln1273_42_fu_12220_p1;

assign grp_fu_21690_p1 = 29'd123;

assign grp_fu_21702_p0 = sext_ln1273_41_fu_12216_p1;

assign grp_fu_21702_p1 = 34'd3741;

assign grp_fu_21714_p0 = sext_ln1273_47_fu_12236_p1;

assign grp_fu_21714_p1 = 35'd5290;

assign grp_fu_21721_p0 = sext_ln1273_40_fu_12212_p1;

assign grp_fu_21721_p1 = 30'd177;

assign grp_fu_21733_p0 = sext_ln1273_45_fu_12232_p1;

assign grp_fu_21733_p1 = 29'd123;

assign grp_fu_21740_p0 = sext_ln1273_44_fu_12228_p1;

assign grp_fu_21740_p1 = 35'd34359733078;

assign grp_fu_21752_p0 = sext_ln1273_42_fu_12220_p1;

assign grp_fu_21752_p1 = 29'd536870789;

assign grp_fu_21764_p0 = sext_ln1273_41_fu_12216_p1;

assign grp_fu_21764_p1 = 34'd17179865443;

assign grp_fu_21776_p0 = sext_ln1273_47_fu_12236_p1;

assign grp_fu_21776_p1 = 35'd34359733078;

assign grp_fu_21783_p0 = sext_ln1273_40_fu_12212_p1;

assign grp_fu_21783_p1 = 30'd1073741647;

assign grp_fu_21795_p0 = sext_ln1273_45_fu_12232_p1;

assign grp_fu_21795_p1 = 29'd536870789;

assign grp_fu_21802_p0 = sext_ln1273_47_reg_23419;

assign grp_fu_21802_p1 = 35'd7479;

assign grp_fu_21810_p0 = sext_ln1273_46_fu_12537_p1;

assign grp_fu_21810_p1 = 28'd47;

assign grp_fu_21819_p0 = sext_ln1273_49_fu_12544_p1;

assign grp_fu_21819_p1 = 35'd7479;

assign grp_fu_21826_p0 = sext_ln1273_48_fu_12540_p1;

assign grp_fu_21826_p1 = 28'd47;

assign grp_fu_21833_p0 = sext_ln1273_44_reg_23405;

assign grp_fu_21833_p1 = 35'd34359730889;

assign grp_fu_21844_p0 = sext_ln1273_43_reg_23399;

assign grp_fu_21844_p1 = 28'd268435409;

assign grp_fu_21855_p0 = sext_ln1273_47_reg_23419;

assign grp_fu_21855_p1 = 35'd34359730889;

assign grp_fu_21863_p0 = sext_ln1273_46_fu_12537_p1;

assign grp_fu_21863_p1 = 28'd268435409;

assign grp_fu_21872_p0 = sext_ln1273_49_fu_12544_p1;

assign grp_fu_21872_p1 = 35'd34359730889;

assign grp_fu_21879_p0 = sext_ln1273_48_fu_12540_p1;

assign grp_fu_21879_p1 = 28'd268435409;

assign grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start = grp_vsub_18_ap_fixed_21_7_0_0_0_s_fu_1177_ap_start_reg;

assign i_2_fu_1298_p2 = (ap_sig_allocacmp_i_1 + 5'd1);

assign icmp_ln74_fu_1292_p2 = ((ap_sig_allocacmp_i_1 == 5'd20) ? 1'b1 : 1'b0);

assign or_ln346_10_fu_8977_p2 = (and_ln896_10_fu_8971_p2 | and_ln895_45_fu_8947_p2);

assign or_ln346_11_fu_9486_p2 = (and_ln896_11_fu_9480_p2 | and_ln895_46_fu_9456_p2);

assign or_ln346_12_fu_9847_p2 = (and_ln896_12_fu_9841_p2 | and_ln895_47_fu_9817_p2);

assign or_ln346_13_fu_10158_p2 = (and_ln896_13_fu_10152_p2 | and_ln895_50_fu_10128_p2);

assign or_ln346_14_fu_2716_p2 = (and_ln896_14_fu_2710_p2 | and_ln895_53_fu_2686_p2);

assign or_ln346_15_fu_4053_p2 = (and_ln896_15_fu_4048_p2 | and_ln895_54_reg_22584);

assign or_ln346_16_fu_4259_p2 = (and_ln896_16_fu_4253_p2 | and_ln895_55_fu_4229_p2);

assign or_ln346_17_fu_5118_p2 = (and_ln896_17_fu_5112_p2 | and_ln895_56_fu_5088_p2);

assign or_ln346_18_fu_6210_p2 = (and_ln896_18_fu_6205_p2 | and_ln895_59_reg_22813);

assign or_ln346_19_fu_6420_p2 = (and_ln896_19_fu_6414_p2 | and_ln895_60_fu_6390_p2);

assign or_ln346_1_fu_2508_p2 = (and_ln896_1_fu_2502_p2 | and_ln895_36_fu_2478_p2);

assign or_ln346_20_fu_7087_p2 = (and_ln896_20_fu_7081_p2 | and_ln895_61_fu_7057_p2);

assign or_ln346_21_fu_7821_p2 = (and_ln896_21_fu_7815_p2 | and_ln895_62_fu_7791_p2);

assign or_ln346_22_fu_8610_p2 = (and_ln896_22_fu_8604_p2 | and_ln895_64_fu_8580_p2);

assign or_ln346_23_fu_9290_p2 = (and_ln896_23_fu_9284_p2 | and_ln895_67_fu_9260_p2);

assign or_ln346_24_fu_2909_p2 = (and_ln896_24_fu_2903_p2 | and_ln895_69_fu_2879_p2);

assign or_ln346_25_fu_4295_p2 = (and_ln896_25_fu_4283_p2 | and_ln895_70_reg_22620);

assign or_ln346_26_fu_6452_p2 = (and_ln896_26_fu_6447_p2 | and_ln895_75_reg_22865);

assign or_ln346_27_fu_6662_p2 = (and_ln896_27_fu_6656_p2 | and_ln895_76_fu_6632_p2);

assign or_ln346_28_fu_7860_p2 = (and_ln896_28_fu_7848_p2 | and_ln895_79_reg_22992);

assign or_ln346_29_fu_8642_p2 = (and_ln896_29_fu_8630_p2 | and_ln895_82_reg_23058);

assign or_ln346_2_fu_3257_p2 = (and_ln896_2_fu_3251_p2 | and_ln895_37_fu_3227_p2);

assign or_ln346_30_fu_10534_p2 = (and_ln896_30_fu_10528_p2 | and_ln895_86_fu_10504_p2);

assign or_ln346_31_fu_11097_p2 = (and_ln896_31_fu_11091_p2 | and_ln895_87_fu_11067_p2);

assign or_ln346_32_fu_11772_p2 = (and_ln896_32_fu_11766_p2 | and_ln895_88_fu_11742_p2);

assign or_ln346_33_fu_10724_p2 = (and_ln896_33_fu_10718_p2 | and_ln895_89_fu_10694_p2);

assign or_ln346_34_fu_11327_p2 = (and_ln896_34_fu_11321_p2 | and_ln895_90_fu_11297_p2);

assign or_ln346_35_fu_11968_p2 = (and_ln896_35_fu_11962_p2 | and_ln895_91_fu_11938_p2);

assign or_ln346_36_fu_10898_p2 = (and_ln896_36_fu_10892_p2 | and_ln895_92_fu_10868_p2);

assign or_ln346_37_fu_11576_p2 = (and_ln896_37_fu_11570_p2 | and_ln895_93_fu_11546_p2);

assign or_ln346_38_fu_12174_p2 = (and_ln896_38_fu_12168_p2 | and_ln895_94_fu_12144_p2);

assign or_ln346_39_fu_13275_p2 = (and_ln896_39_fu_13269_p2 | and_ln895_95_fu_13245_p2);

assign or_ln346_3_fu_4010_p2 = (and_ln896_3_fu_4004_p2 | and_ln895_38_fu_3980_p2);

assign or_ln346_40_fu_13449_p2 = (and_ln896_40_fu_13443_p2 | and_ln895_98_fu_13419_p2);

assign or_ln346_41_fu_13619_p2 = (and_ln896_41_fu_13613_p2 | and_ln895_101_fu_13589_p2);

assign or_ln346_42_fu_17161_p2 = (and_ln896_42_fu_17149_p2 | and_ln895_102_reg_23629);

assign or_ln346_43_fu_13809_p2 = (and_ln896_43_fu_13803_p2 | and_ln895_104_fu_13779_p2);

assign or_ln346_44_fu_17249_p2 = (and_ln896_44_fu_17237_p2 | and_ln895_105_reg_23665);

assign or_ln346_45_fu_13983_p2 = (and_ln896_45_fu_13977_p2 | and_ln895_107_fu_13953_p2);

assign or_ln346_46_fu_15711_p2 = (and_ln896_46_fu_15705_p2 | and_ln895_108_fu_15681_p2);

assign or_ln346_47_fu_17505_p2 = (and_ln896_47_fu_17491_p2 | and_ln895_109_fu_17467_p2);

assign or_ln346_48_fu_14180_p2 = (and_ln896_48_fu_14174_p2 | and_ln895_110_fu_14150_p2);

assign or_ln346_49_fu_15948_p2 = (and_ln896_49_fu_15942_p2 | and_ln895_111_fu_15918_p2);

assign or_ln346_4_fu_4851_p2 = (and_ln896_4_fu_4845_p2 | and_ln895_39_fu_4821_p2);

assign or_ln346_50_fu_17717_p2 = (and_ln896_50_fu_17703_p2 | and_ln895_112_fu_17679_p2);

assign or_ln346_51_fu_16141_p2 = (and_ln896_51_fu_16135_p2 | and_ln895_113_fu_16111_p2);

assign or_ln346_52_fu_16315_p2 = (and_ln896_52_fu_16309_p2 | and_ln895_116_fu_16285_p2);

assign or_ln346_53_fu_14357_p2 = (and_ln896_53_fu_14351_p2 | and_ln895_119_fu_14327_p2);

assign or_ln346_54_fu_17989_p2 = (and_ln896_54_fu_17977_p2 | and_ln895_120_reg_23763);

assign or_ln346_55_fu_14547_p2 = (and_ln896_55_fu_14541_p2 | and_ln895_122_fu_14517_p2);

assign or_ln346_56_fu_18077_p2 = (and_ln896_56_fu_18065_p2 | and_ln895_123_reg_23799);

assign or_ln346_57_fu_14721_p2 = (and_ln896_57_fu_14715_p2 | and_ln895_125_fu_14691_p2);

assign or_ln346_58_fu_16869_p2 = (and_ln896_58_fu_16863_p2 | and_ln895_126_fu_16839_p2);

assign or_ln346_59_fu_18333_p2 = (and_ln896_59_fu_18319_p2 | and_ln895_127_fu_18295_p2);

assign or_ln346_5_fu_5472_p2 = (and_ln896_5_fu_5466_p2 | and_ln895_40_fu_5442_p2);

assign or_ln346_60_fu_14918_p2 = (and_ln896_60_fu_14912_p2 | and_ln895_128_fu_14888_p2);

assign or_ln346_61_fu_17106_p2 = (and_ln896_61_fu_17100_p2 | and_ln895_129_fu_17076_p2);

assign or_ln346_62_fu_18545_p2 = (and_ln896_62_fu_18531_p2 | and_ln895_130_fu_18507_p2);

assign or_ln346_63_fu_12459_p2 = (and_ln896_64_fu_12445_p2 | and_ln895_134_fu_12427_p2);

assign or_ln346_64_fu_12616_p2 = (and_ln896_66_fu_12602_p2 | and_ln895_136_fu_12584_p2);

assign or_ln346_65_fu_12726_p2 = (and_ln896_68_fu_12712_p2 | and_ln895_137_fu_12694_p2);

assign or_ln346_66_fu_12947_p2 = (and_ln896_70_fu_12933_p2 | and_ln895_140_fu_12915_p2);

assign or_ln346_67_fu_13096_p2 = (and_ln896_72_fu_13082_p2 | and_ln895_142_fu_13064_p2);

assign or_ln346_6_fu_6162_p2 = (and_ln896_6_fu_6156_p2 | and_ln895_41_fu_6132_p2);

assign or_ln346_7_fu_6858_p2 = (and_ln896_7_fu_6852_p2 | and_ln895_42_fu_6828_p2);

assign or_ln346_8_fu_7570_p2 = (and_ln896_8_fu_7564_p2 | and_ln895_43_fu_7540_p2);

assign or_ln346_9_fu_8363_p2 = (and_ln896_9_fu_8357_p2 | and_ln895_44_fu_8333_p2);

assign or_ln346_fu_2141_p2 = (and_ln896_fu_2135_p2 | and_ln895_35_fu_2111_p2);

assign or_ln888_10_fu_8885_p2 = (xor_ln888_20_fu_8879_p2 | tmp_134_fu_8851_p3);

assign or_ln888_11_fu_9394_p2 = (xor_ln888_22_fu_9388_p2 | tmp_140_fu_9360_p3);

assign or_ln888_12_fu_9755_p2 = (xor_ln888_24_fu_9749_p2 | tmp_146_fu_9721_p3);

assign or_ln888_13_fu_10066_p2 = (xor_ln888_26_fu_10060_p2 | tmp_156_fu_10032_p3);

assign or_ln888_14_fu_2625_p2 = (xor_ln888_28_fu_2619_p2 | tmp_166_fu_2592_p3);

assign or_ln888_15_fu_3402_p2 = (xor_ln888_30_fu_3396_p2 | tmp_172_fu_3374_p3);

assign or_ln888_16_fu_4167_p2 = (xor_ln888_32_fu_4161_p2 | tmp_178_fu_4133_p3);

assign or_ln888_17_fu_5026_p2 = (xor_ln888_34_fu_5020_p2 | tmp_184_fu_4992_p3);

assign or_ln888_18_fu_5710_p2 = (xor_ln888_36_fu_5704_p2 | tmp_194_fu_5682_p3);

assign or_ln888_19_fu_6328_p2 = (xor_ln888_38_fu_6322_p2 | tmp_200_fu_6294_p3);

assign or_ln888_1_fu_2416_p2 = (xor_ln888_2_fu_2410_p2 | tmp_80_fu_2382_p3);

assign or_ln888_20_fu_6995_p2 = (xor_ln888_40_fu_6989_p2 | tmp_206_fu_6961_p3);

assign or_ln888_21_fu_7729_p2 = (xor_ln888_42_fu_7723_p2 | tmp_212_fu_7695_p3);

assign or_ln888_22_fu_8518_p2 = (xor_ln888_44_fu_8512_p2 | tmp_220_fu_8484_p3);

assign or_ln888_23_fu_9198_p2 = (xor_ln888_46_fu_9192_p2 | tmp_230_fu_9164_p3);

assign or_ln888_24_fu_2818_p2 = (xor_ln888_48_fu_2812_p2 | tmp_238_fu_2785_p3);

assign or_ln888_25_fu_3576_p2 = (xor_ln888_50_fu_3570_p2 | tmp_244_fu_3548_p3);

assign or_ln888_26_fu_5891_p2 = (xor_ln888_52_fu_5885_p2 | tmp_258_fu_5863_p3);

assign or_ln888_27_fu_6570_p2 = (xor_ln888_54_fu_6564_p2 | tmp_264_fu_6536_p3);

assign or_ln888_28_fu_7310_p2 = (xor_ln888_56_fu_7304_p2 | tmp_274_fu_7282_p3);

assign or_ln888_29_fu_8060_p2 = (xor_ln888_58_fu_8054_p2 | tmp_284_fu_8032_p3);

assign or_ln888_2_fu_3165_p2 = (xor_ln888_4_fu_3159_p2 | tmp_86_fu_3131_p3);

assign or_ln888_30_fu_10443_p2 = (xor_ln888_60_fu_10437_p2 | tmp_296_fu_10410_p3);

assign or_ln888_31_fu_11005_p2 = (xor_ln888_62_fu_10999_p2 | tmp_302_fu_10971_p3);

assign or_ln888_32_fu_11680_p2 = (xor_ln888_64_fu_11674_p2 | tmp_308_fu_11646_p3);

assign or_ln888_33_fu_10633_p2 = (xor_ln888_66_fu_10627_p2 | tmp_314_fu_10600_p3);

assign or_ln888_34_fu_11235_p2 = (xor_ln888_68_fu_11229_p2 | tmp_320_fu_11201_p3);

assign or_ln888_35_fu_11876_p2 = (xor_ln888_70_fu_11870_p2 | tmp_326_fu_11842_p3);

assign or_ln888_36_fu_10807_p2 = (xor_ln888_72_fu_10801_p2 | tmp_332_fu_10774_p3);

assign or_ln888_37_fu_11484_p2 = (xor_ln888_74_fu_11478_p2 | tmp_338_fu_11450_p3);

assign or_ln888_38_fu_12082_p2 = (xor_ln888_76_fu_12076_p2 | tmp_344_fu_12048_p3);

assign or_ln888_39_fu_13184_p2 = (xor_ln888_78_fu_13178_p2 | tmp_350_fu_13151_p3);

assign or_ln888_3_fu_3918_p2 = (xor_ln888_6_fu_3912_p2 | tmp_92_fu_3884_p3);

assign or_ln888_40_fu_13358_p2 = (xor_ln888_80_fu_13352_p2 | tmp_360_fu_13325_p3);

assign or_ln888_41_fu_13528_p2 = (xor_ln888_82_fu_13522_p2 | tmp_370_fu_13495_p3);

assign or_ln888_42_fu_15259_p2 = (xor_ln888_84_fu_15253_p2 | tmp_376_fu_15231_p3);

assign or_ln888_43_fu_13718_p2 = (xor_ln888_86_fu_13712_p2 | tmp_384_fu_13685_p3);

assign or_ln888_44_fu_15451_p2 = (xor_ln888_88_fu_15445_p2 | tmp_390_fu_15423_p3);

assign or_ln888_45_fu_13892_p2 = (xor_ln888_90_fu_13886_p2 | tmp_398_fu_13859_p3);

assign or_ln888_46_fu_15619_p2 = (xor_ln888_92_fu_15613_p2 | tmp_404_fu_15585_p3);

assign or_ln888_47_fu_17405_p2 = (xor_ln888_94_fu_17399_p2 | tmp_410_fu_17371_p3);

assign or_ln888_48_fu_14089_p2 = (xor_ln888_96_fu_14083_p2 | tmp_416_fu_14056_p3);

assign or_ln888_49_fu_15856_p2 = (xor_ln888_98_fu_15850_p2 | tmp_422_fu_15822_p3);

assign or_ln888_4_fu_4759_p2 = (xor_ln888_8_fu_4753_p2 | tmp_98_fu_4725_p3);

assign or_ln888_50_fu_17617_p2 = (xor_ln888_100_fu_17611_p2 | tmp_428_fu_17583_p3);

assign or_ln888_51_fu_16050_p2 = (xor_ln888_102_fu_16044_p2 | tmp_434_fu_16017_p3);

assign or_ln888_52_fu_16224_p2 = (xor_ln888_104_fu_16218_p2 | tmp_444_fu_16191_p3);

assign or_ln888_53_fu_14266_p2 = (xor_ln888_106_fu_14260_p2 | tmp_454_fu_14233_p3);

assign or_ln888_54_fu_16417_p2 = (xor_ln888_108_fu_16411_p2 | tmp_460_fu_16389_p3);

assign or_ln888_55_fu_14456_p2 = (xor_ln888_110_fu_14450_p2 | tmp_468_fu_14423_p3);

assign or_ln888_56_fu_16609_p2 = (xor_ln888_112_fu_16603_p2 | tmp_474_fu_16581_p3);

assign or_ln888_57_fu_14630_p2 = (xor_ln888_114_fu_14624_p2 | tmp_482_fu_14597_p3);

assign or_ln888_58_fu_16777_p2 = (xor_ln888_116_fu_16771_p2 | tmp_488_fu_16743_p3);

assign or_ln888_59_fu_18233_p2 = (xor_ln888_118_fu_18227_p2 | tmp_494_fu_18199_p3);

assign or_ln888_5_fu_5380_p2 = (xor_ln888_10_fu_5374_p2 | tmp_104_fu_5346_p3);

assign or_ln888_60_fu_14827_p2 = (xor_ln888_120_fu_14821_p2 | tmp_500_fu_14794_p3);

assign or_ln888_61_fu_17014_p2 = (xor_ln888_122_fu_17008_p2 | tmp_506_fu_16980_p3);

assign or_ln888_62_fu_18445_p2 = (xor_ln888_124_fu_18439_p2 | tmp_512_fu_18411_p3);

assign or_ln888_6_fu_6070_p2 = (xor_ln888_12_fu_6064_p2 | tmp_110_fu_6036_p3);

assign or_ln888_7_fu_6766_p2 = (xor_ln888_14_fu_6760_p2 | tmp_116_fu_6732_p3);

assign or_ln888_8_fu_7478_p2 = (xor_ln888_16_fu_7472_p2 | tmp_122_fu_7444_p3);

assign or_ln888_9_fu_8271_p2 = (xor_ln888_18_fu_8265_p2 | tmp_128_fu_8237_p3);

assign or_ln888_fu_2050_p2 = (xor_ln888_fu_2044_p2 | tmp_74_fu_2017_p3);

assign or_ln890_10_fu_8911_p2 = (xor_ln890_10_fu_8905_p2 | or_ln888_10_fu_8885_p2);

assign or_ln890_11_fu_9420_p2 = (xor_ln890_11_fu_9414_p2 | or_ln888_11_fu_9394_p2);

assign or_ln890_12_fu_9781_p2 = (xor_ln890_12_fu_9775_p2 | or_ln888_12_fu_9755_p2);

assign or_ln890_13_fu_10092_p2 = (xor_ln890_13_fu_10086_p2 | or_ln888_13_fu_10066_p2);

assign or_ln890_14_fu_2650_p2 = (xor_ln890_14_fu_2644_p2 | or_ln888_14_fu_2625_p2);

assign or_ln890_15_fu_3428_p2 = (xor_ln890_15_fu_3422_p2 | or_ln888_15_fu_3402_p2);

assign or_ln890_16_fu_4193_p2 = (xor_ln890_16_fu_4187_p2 | or_ln888_16_fu_4167_p2);

assign or_ln890_17_fu_5052_p2 = (xor_ln890_17_fu_5046_p2 | or_ln888_17_fu_5026_p2);

assign or_ln890_18_fu_5736_p2 = (xor_ln890_18_fu_5730_p2 | or_ln888_18_fu_5710_p2);

assign or_ln890_19_fu_6354_p2 = (xor_ln890_19_fu_6348_p2 | or_ln888_19_fu_6328_p2);

assign or_ln890_1_fu_2442_p2 = (xor_ln890_1_fu_2436_p2 | or_ln888_1_fu_2416_p2);

assign or_ln890_20_fu_7021_p2 = (xor_ln890_20_fu_7015_p2 | or_ln888_20_fu_6995_p2);

assign or_ln890_21_fu_7755_p2 = (xor_ln890_21_fu_7749_p2 | or_ln888_21_fu_7729_p2);

assign or_ln890_22_fu_8544_p2 = (xor_ln890_22_fu_8538_p2 | or_ln888_22_fu_8518_p2);

assign or_ln890_23_fu_9224_p2 = (xor_ln890_23_fu_9218_p2 | or_ln888_23_fu_9198_p2);

assign or_ln890_24_fu_2843_p2 = (xor_ln890_24_fu_2837_p2 | or_ln888_24_fu_2818_p2);

assign or_ln890_25_fu_3602_p2 = (xor_ln890_25_fu_3596_p2 | or_ln888_25_fu_3576_p2);

assign or_ln890_26_fu_5917_p2 = (xor_ln890_26_fu_5911_p2 | or_ln888_26_fu_5891_p2);

assign or_ln890_27_fu_6596_p2 = (xor_ln890_27_fu_6590_p2 | or_ln888_27_fu_6570_p2);

assign or_ln890_28_fu_7336_p2 = (xor_ln890_28_fu_7330_p2 | or_ln888_28_fu_7310_p2);

assign or_ln890_29_fu_8086_p2 = (xor_ln890_29_fu_8080_p2 | or_ln888_29_fu_8060_p2);

assign or_ln890_2_fu_3191_p2 = (xor_ln890_2_fu_3185_p2 | or_ln888_2_fu_3165_p2);

assign or_ln890_30_fu_10468_p2 = (xor_ln890_30_fu_10462_p2 | or_ln888_30_fu_10443_p2);

assign or_ln890_31_fu_11031_p2 = (xor_ln890_31_fu_11025_p2 | or_ln888_31_fu_11005_p2);

assign or_ln890_32_fu_11706_p2 = (xor_ln890_32_fu_11700_p2 | or_ln888_32_fu_11680_p2);

assign or_ln890_33_fu_10658_p2 = (xor_ln890_33_fu_10652_p2 | or_ln888_33_fu_10633_p2);

assign or_ln890_34_fu_11261_p2 = (xor_ln890_34_fu_11255_p2 | or_ln888_34_fu_11235_p2);

assign or_ln890_35_fu_11902_p2 = (xor_ln890_35_fu_11896_p2 | or_ln888_35_fu_11876_p2);

assign or_ln890_36_fu_10832_p2 = (xor_ln890_36_fu_10826_p2 | or_ln888_36_fu_10807_p2);

assign or_ln890_37_fu_11510_p2 = (xor_ln890_37_fu_11504_p2 | or_ln888_37_fu_11484_p2);

assign or_ln890_38_fu_12108_p2 = (xor_ln890_38_fu_12102_p2 | or_ln888_38_fu_12082_p2);

assign or_ln890_39_fu_13209_p2 = (xor_ln890_39_fu_13203_p2 | or_ln888_39_fu_13184_p2);

assign or_ln890_3_fu_3944_p2 = (xor_ln890_3_fu_3938_p2 | or_ln888_3_fu_3918_p2);

assign or_ln890_40_fu_13383_p2 = (xor_ln890_40_fu_13377_p2 | or_ln888_40_fu_13358_p2);

assign or_ln890_41_fu_13553_p2 = (xor_ln890_41_fu_13547_p2 | or_ln888_41_fu_13528_p2);

assign or_ln890_42_fu_15285_p2 = (xor_ln890_42_fu_15279_p2 | or_ln888_42_fu_15259_p2);

assign or_ln890_43_fu_13743_p2 = (xor_ln890_43_fu_13737_p2 | or_ln888_43_fu_13718_p2);

assign or_ln890_44_fu_15477_p2 = (xor_ln890_44_fu_15471_p2 | or_ln888_44_fu_15451_p2);

assign or_ln890_45_fu_13917_p2 = (xor_ln890_45_fu_13911_p2 | or_ln888_45_fu_13892_p2);

assign or_ln890_46_fu_15645_p2 = (xor_ln890_46_fu_15639_p2 | or_ln888_46_fu_15619_p2);

assign or_ln890_47_fu_17431_p2 = (xor_ln890_47_fu_17425_p2 | or_ln888_47_fu_17405_p2);

assign or_ln890_48_fu_14114_p2 = (xor_ln890_48_fu_14108_p2 | or_ln888_48_fu_14089_p2);

assign or_ln890_49_fu_15882_p2 = (xor_ln890_49_fu_15876_p2 | or_ln888_49_fu_15856_p2);

assign or_ln890_4_fu_4785_p2 = (xor_ln890_4_fu_4779_p2 | or_ln888_4_fu_4759_p2);

assign or_ln890_50_fu_17643_p2 = (xor_ln890_50_fu_17637_p2 | or_ln888_50_fu_17617_p2);

assign or_ln890_51_fu_16075_p2 = (xor_ln890_51_fu_16069_p2 | or_ln888_51_fu_16050_p2);

assign or_ln890_52_fu_16249_p2 = (xor_ln890_52_fu_16243_p2 | or_ln888_52_fu_16224_p2);

assign or_ln890_53_fu_14291_p2 = (xor_ln890_53_fu_14285_p2 | or_ln888_53_fu_14266_p2);

assign or_ln890_54_fu_16443_p2 = (xor_ln890_54_fu_16437_p2 | or_ln888_54_fu_16417_p2);

assign or_ln890_55_fu_14481_p2 = (xor_ln890_55_fu_14475_p2 | or_ln888_55_fu_14456_p2);

assign or_ln890_56_fu_16635_p2 = (xor_ln890_56_fu_16629_p2 | or_ln888_56_fu_16609_p2);

assign or_ln890_57_fu_14655_p2 = (xor_ln890_57_fu_14649_p2 | or_ln888_57_fu_14630_p2);

assign or_ln890_58_fu_16803_p2 = (xor_ln890_58_fu_16797_p2 | or_ln888_58_fu_16777_p2);

assign or_ln890_59_fu_18259_p2 = (xor_ln890_59_fu_18253_p2 | or_ln888_59_fu_18233_p2);

assign or_ln890_5_fu_5406_p2 = (xor_ln890_5_fu_5400_p2 | or_ln888_5_fu_5380_p2);

assign or_ln890_60_fu_14852_p2 = (xor_ln890_60_fu_14846_p2 | or_ln888_60_fu_14827_p2);

assign or_ln890_61_fu_17040_p2 = (xor_ln890_61_fu_17034_p2 | or_ln888_61_fu_17014_p2);

assign or_ln890_62_fu_18471_p2 = (xor_ln890_62_fu_18465_p2 | or_ln888_62_fu_18445_p2);

assign or_ln890_6_fu_6096_p2 = (xor_ln890_6_fu_6090_p2 | or_ln888_6_fu_6070_p2);

assign or_ln890_7_fu_6792_p2 = (xor_ln890_7_fu_6786_p2 | or_ln888_7_fu_6766_p2);

assign or_ln890_8_fu_7504_p2 = (xor_ln890_8_fu_7498_p2 | or_ln888_8_fu_7478_p2);

assign or_ln890_9_fu_8297_p2 = (xor_ln890_9_fu_8291_p2 | or_ln888_9_fu_8271_p2);

assign or_ln890_fu_2075_p2 = (xor_ln890_fu_2069_p2 | or_ln888_fu_2050_p2);

assign or_ln895_10_fu_8935_p2 = (xor_ln895_47_fu_8929_p2 | tmp_134_fu_8851_p3);

assign or_ln895_11_fu_9444_p2 = (xor_ln895_49_fu_9438_p2 | tmp_140_fu_9360_p3);

assign or_ln895_12_fu_9805_p2 = (xor_ln895_51_fu_9799_p2 | tmp_146_fu_9721_p3);

assign or_ln895_13_fu_10116_p2 = (xor_ln895_55_fu_10110_p2 | tmp_156_fu_10032_p3);

assign or_ln895_14_fu_2674_p2 = (xor_ln895_59_fu_2668_p2 | tmp_166_fu_2592_p3);

assign or_ln895_15_fu_3446_p2 = (xor_ln895_61_fu_3440_p2 | tmp_172_fu_3374_p3);

assign or_ln895_16_fu_4217_p2 = (xor_ln895_63_fu_4211_p2 | tmp_178_fu_4133_p3);

assign or_ln895_17_fu_5076_p2 = (xor_ln895_65_fu_5070_p2 | tmp_184_fu_4992_p3);

assign or_ln895_18_fu_5754_p2 = (xor_ln895_69_fu_5748_p2 | tmp_194_fu_5682_p3);

assign or_ln895_19_fu_6378_p2 = (xor_ln895_71_fu_6372_p2 | tmp_200_fu_6294_p3);

assign or_ln895_1_fu_2466_p2 = (xor_ln895_29_fu_2460_p2 | tmp_80_fu_2382_p3);

assign or_ln895_20_fu_7045_p2 = (xor_ln895_73_fu_7039_p2 | tmp_206_fu_6961_p3);

assign or_ln895_21_fu_7779_p2 = (xor_ln895_75_fu_7773_p2 | tmp_212_fu_7695_p3);

assign or_ln895_22_fu_8568_p2 = (xor_ln895_78_fu_8562_p2 | tmp_220_fu_8484_p3);

assign or_ln895_23_fu_9248_p2 = (xor_ln895_82_fu_9242_p2 | tmp_230_fu_9164_p3);

assign or_ln895_24_fu_2867_p2 = (xor_ln895_85_fu_2861_p2 | tmp_238_fu_2785_p3);

assign or_ln895_25_fu_3620_p2 = (xor_ln895_87_fu_3614_p2 | tmp_244_fu_3548_p3);

assign or_ln895_26_fu_5935_p2 = (xor_ln895_93_fu_5929_p2 | tmp_258_fu_5863_p3);

assign or_ln895_27_fu_6620_p2 = (xor_ln895_95_fu_6614_p2 | tmp_264_fu_6536_p3);

assign or_ln895_28_fu_7354_p2 = (xor_ln895_99_fu_7348_p2 | tmp_274_fu_7282_p3);

assign or_ln895_29_fu_8104_p2 = (xor_ln895_103_fu_8098_p2 | tmp_284_fu_8032_p3);

assign or_ln895_2_fu_3215_p2 = (xor_ln895_31_fu_3209_p2 | tmp_86_fu_3131_p3);

assign or_ln895_30_fu_10492_p2 = (xor_ln895_108_fu_10486_p2 | tmp_296_fu_10410_p3);

assign or_ln895_31_fu_11055_p2 = (xor_ln895_110_fu_11049_p2 | tmp_302_fu_10971_p3);

assign or_ln895_32_fu_11730_p2 = (xor_ln895_112_fu_11724_p2 | tmp_308_fu_11646_p3);

assign or_ln895_33_fu_10682_p2 = (xor_ln895_114_fu_10676_p2 | tmp_314_fu_10600_p3);

assign or_ln895_34_fu_11285_p2 = (xor_ln895_116_fu_11279_p2 | tmp_320_fu_11201_p3);

assign or_ln895_35_fu_11926_p2 = (xor_ln895_118_fu_11920_p2 | tmp_326_fu_11842_p3);

assign or_ln895_36_fu_10856_p2 = (xor_ln895_120_fu_10850_p2 | tmp_332_fu_10774_p3);

assign or_ln895_37_fu_11534_p2 = (xor_ln895_122_fu_11528_p2 | tmp_338_fu_11450_p3);

assign or_ln895_38_fu_12132_p2 = (xor_ln895_124_fu_12126_p2 | tmp_344_fu_12048_p3);

assign or_ln895_39_fu_13233_p2 = (xor_ln895_126_fu_13227_p2 | tmp_350_fu_13151_p3);

assign or_ln895_3_fu_3968_p2 = (xor_ln895_33_fu_3962_p2 | tmp_92_fu_3884_p3);

assign or_ln895_40_fu_13407_p2 = (xor_ln895_130_fu_13401_p2 | tmp_360_fu_13325_p3);

assign or_ln895_41_fu_13577_p2 = (xor_ln895_134_fu_13571_p2 | tmp_370_fu_13495_p3);

assign or_ln895_42_fu_15303_p2 = (xor_ln895_136_fu_15297_p2 | tmp_376_fu_15231_p3);

assign or_ln895_43_fu_13767_p2 = (xor_ln895_139_fu_13761_p2 | tmp_384_fu_13685_p3);

assign or_ln895_44_fu_15495_p2 = (xor_ln895_141_fu_15489_p2 | tmp_390_fu_15423_p3);

assign or_ln895_45_fu_13941_p2 = (xor_ln895_144_fu_13935_p2 | tmp_398_fu_13859_p3);

assign or_ln895_46_fu_15669_p2 = (xor_ln895_146_fu_15663_p2 | tmp_404_fu_15585_p3);

assign or_ln895_47_fu_17455_p2 = (xor_ln895_148_fu_17449_p2 | tmp_410_fu_17371_p3);

assign or_ln895_48_fu_14138_p2 = (xor_ln895_150_fu_14132_p2 | tmp_416_fu_14056_p3);

assign or_ln895_49_fu_15906_p2 = (xor_ln895_152_fu_15900_p2 | tmp_422_fu_15822_p3);

assign or_ln895_4_fu_4809_p2 = (xor_ln895_35_fu_4803_p2 | tmp_98_fu_4725_p3);

assign or_ln895_50_fu_17667_p2 = (xor_ln895_154_fu_17661_p2 | tmp_428_fu_17583_p3);

assign or_ln895_51_fu_16099_p2 = (xor_ln895_156_fu_16093_p2 | tmp_434_fu_16017_p3);

assign or_ln895_52_fu_16273_p2 = (xor_ln895_160_fu_16267_p2 | tmp_444_fu_16191_p3);

assign or_ln895_53_fu_14315_p2 = (xor_ln895_164_fu_14309_p2 | tmp_454_fu_14233_p3);

assign or_ln895_54_fu_16461_p2 = (xor_ln895_166_fu_16455_p2 | tmp_460_fu_16389_p3);

assign or_ln895_55_fu_14505_p2 = (xor_ln895_169_fu_14499_p2 | tmp_468_fu_14423_p3);

assign or_ln895_56_fu_16653_p2 = (xor_ln895_171_fu_16647_p2 | tmp_474_fu_16581_p3);

assign or_ln895_57_fu_14679_p2 = (xor_ln895_174_fu_14673_p2 | tmp_482_fu_14597_p3);

assign or_ln895_58_fu_16827_p2 = (xor_ln895_176_fu_16821_p2 | tmp_488_fu_16743_p3);

assign or_ln895_59_fu_18283_p2 = (xor_ln895_178_fu_18277_p2 | tmp_494_fu_18199_p3);

assign or_ln895_5_fu_5430_p2 = (xor_ln895_37_fu_5424_p2 | tmp_104_fu_5346_p3);

assign or_ln895_60_fu_14876_p2 = (xor_ln895_180_fu_14870_p2 | tmp_500_fu_14794_p3);

assign or_ln895_61_fu_17064_p2 = (xor_ln895_182_fu_17058_p2 | tmp_506_fu_16980_p3);

assign or_ln895_62_fu_18495_p2 = (xor_ln895_184_fu_18489_p2 | tmp_512_fu_18411_p3);

assign or_ln895_63_fu_12415_p2 = (tmp_523_fu_12407_p3 | tmp_522_fu_12399_p3);

assign or_ln895_64_fu_12572_p2 = (tmp_528_fu_12564_p3 | tmp_527_fu_12556_p3);

assign or_ln895_65_fu_12682_p2 = (tmp_531_fu_12674_p3 | tmp_530_fu_12666_p3);

assign or_ln895_66_fu_12903_p2 = (tmp_538_fu_12895_p3 | tmp_537_fu_12887_p3);

assign or_ln895_67_fu_13052_p2 = (tmp_543_fu_13044_p3 | tmp_542_fu_13036_p3);

assign or_ln895_6_fu_6120_p2 = (xor_ln895_39_fu_6114_p2 | tmp_110_fu_6036_p3);

assign or_ln895_7_fu_6816_p2 = (xor_ln895_41_fu_6810_p2 | tmp_116_fu_6732_p3);

assign or_ln895_8_fu_7528_p2 = (xor_ln895_43_fu_7522_p2 | tmp_122_fu_7444_p3);

assign or_ln895_9_fu_8321_p2 = (xor_ln895_45_fu_8315_p2 | tmp_128_fu_8237_p3);

assign or_ln895_fu_2099_p2 = (xor_ln895_27_fu_2093_p2 | tmp_74_fu_2017_p3);

assign or_ln896_10_fu_8959_p2 = (xor_ln896_21_fu_8953_p2 | xor_ln896_20_fu_8859_p2);

assign or_ln896_11_fu_9468_p2 = (xor_ln896_23_fu_9462_p2 | xor_ln896_22_fu_9368_p2);

assign or_ln896_12_fu_9829_p2 = (xor_ln896_25_fu_9823_p2 | xor_ln896_24_fu_9729_p2);

assign or_ln896_13_fu_10140_p2 = (xor_ln896_29_fu_10134_p2 | xor_ln896_28_fu_10040_p2);

assign or_ln896_14_fu_2698_p2 = (xor_ln896_33_fu_2692_p2 | xor_ln896_32_fu_2600_p2);

assign or_ln896_15_fu_3470_p2 = (xor_ln896_35_fu_3464_p2 | xor_ln896_34_fu_3382_p2);

assign or_ln896_16_fu_4241_p2 = (xor_ln896_37_fu_4235_p2 | xor_ln896_36_fu_4141_p2);

assign or_ln896_17_fu_5100_p2 = (xor_ln896_39_fu_5094_p2 | xor_ln896_38_fu_5000_p2);

assign or_ln896_18_fu_5778_p2 = (xor_ln896_43_fu_5772_p2 | xor_ln896_42_fu_5690_p2);

assign or_ln896_19_fu_6402_p2 = (xor_ln896_45_fu_6396_p2 | xor_ln896_44_fu_6302_p2);

assign or_ln896_1_fu_2490_p2 = (xor_ln896_3_fu_2484_p2 | xor_ln896_2_fu_2390_p2);

assign or_ln896_20_fu_7069_p2 = (xor_ln896_47_fu_7063_p2 | xor_ln896_46_fu_6969_p2);

assign or_ln896_21_fu_7803_p2 = (xor_ln896_49_fu_7797_p2 | xor_ln896_48_fu_7703_p2);

assign or_ln896_22_fu_8592_p2 = (xor_ln896_52_fu_8586_p2 | xor_ln896_51_fu_8492_p2);

assign or_ln896_23_fu_9272_p2 = (xor_ln896_56_fu_9266_p2 | xor_ln896_55_fu_9172_p2);

assign or_ln896_24_fu_2891_p2 = (xor_ln896_59_fu_2885_p2 | xor_ln896_58_fu_2793_p2);

assign or_ln896_25_fu_3644_p2 = (xor_ln896_61_fu_3638_p2 | xor_ln896_60_fu_3556_p2);

assign or_ln896_26_fu_5959_p2 = (xor_ln896_67_fu_5953_p2 | xor_ln896_66_fu_5871_p2);

assign or_ln896_27_fu_6644_p2 = (xor_ln896_69_fu_6638_p2 | xor_ln896_68_fu_6544_p2);

assign or_ln896_28_fu_7378_p2 = (xor_ln896_73_fu_7372_p2 | xor_ln896_72_fu_7290_p2);

assign or_ln896_29_fu_8128_p2 = (xor_ln896_77_fu_8122_p2 | xor_ln896_76_fu_8040_p2);

assign or_ln896_2_fu_3239_p2 = (xor_ln896_5_fu_3233_p2 | xor_ln896_4_fu_3139_p2);

assign or_ln896_30_fu_10516_p2 = (xor_ln896_79_fu_10510_p2 | xor_ln896_78_fu_10418_p2);

assign or_ln896_31_fu_11079_p2 = (xor_ln896_81_fu_11073_p2 | xor_ln896_80_fu_10979_p2);

assign or_ln896_32_fu_11754_p2 = (xor_ln896_83_fu_11748_p2 | xor_ln896_82_fu_11654_p2);

assign or_ln896_33_fu_10706_p2 = (xor_ln896_85_fu_10700_p2 | xor_ln896_84_fu_10608_p2);

assign or_ln896_34_fu_11309_p2 = (xor_ln896_87_fu_11303_p2 | xor_ln896_86_fu_11209_p2);

assign or_ln896_35_fu_11950_p2 = (xor_ln896_89_fu_11944_p2 | xor_ln896_88_fu_11850_p2);

assign or_ln896_36_fu_10880_p2 = (xor_ln896_91_fu_10874_p2 | xor_ln896_90_fu_10782_p2);

assign or_ln896_37_fu_11558_p2 = (xor_ln896_93_fu_11552_p2 | xor_ln896_92_fu_11458_p2);

assign or_ln896_38_fu_12156_p2 = (xor_ln896_95_fu_12150_p2 | xor_ln896_94_fu_12056_p2);

assign or_ln896_39_fu_13257_p2 = (xor_ln896_97_fu_13251_p2 | xor_ln896_96_fu_13159_p2);

assign or_ln896_3_fu_3992_p2 = (xor_ln896_7_fu_3986_p2 | xor_ln896_6_fu_3892_p2);

assign or_ln896_40_fu_13431_p2 = (xor_ln896_101_fu_13425_p2 | xor_ln896_100_fu_13333_p2);

assign or_ln896_41_fu_13601_p2 = (xor_ln896_105_fu_13595_p2 | xor_ln896_104_fu_13503_p2);

assign or_ln896_42_fu_15327_p2 = (xor_ln896_107_fu_15321_p2 | xor_ln896_106_fu_15239_p2);

assign or_ln896_43_fu_13791_p2 = (xor_ln896_110_fu_13785_p2 | xor_ln896_109_fu_13693_p2);

assign or_ln896_44_fu_15519_p2 = (xor_ln896_112_fu_15513_p2 | xor_ln896_111_fu_15431_p2);

assign or_ln896_45_fu_13965_p2 = (xor_ln896_115_fu_13959_p2 | xor_ln896_114_fu_13867_p2);

assign or_ln896_46_fu_15693_p2 = (xor_ln896_117_fu_15687_p2 | xor_ln896_116_fu_15593_p2);

assign or_ln896_47_fu_17479_p2 = (xor_ln896_119_fu_17473_p2 | xor_ln896_118_fu_17379_p2);

assign or_ln896_48_fu_14162_p2 = (xor_ln896_121_fu_14156_p2 | xor_ln896_120_fu_14064_p2);

assign or_ln896_49_fu_15930_p2 = (xor_ln896_123_fu_15924_p2 | xor_ln896_122_fu_15830_p2);

assign or_ln896_4_fu_4833_p2 = (xor_ln896_9_fu_4827_p2 | xor_ln896_8_fu_4733_p2);

assign or_ln896_50_fu_17691_p2 = (xor_ln896_125_fu_17685_p2 | xor_ln896_124_fu_17591_p2);

assign or_ln896_51_fu_16123_p2 = (xor_ln896_127_fu_16117_p2 | xor_ln896_126_fu_16025_p2);

assign or_ln896_52_fu_16297_p2 = (xor_ln896_131_fu_16291_p2 | xor_ln896_130_fu_16199_p2);

assign or_ln896_53_fu_14339_p2 = (xor_ln896_135_fu_14333_p2 | xor_ln896_134_fu_14241_p2);

assign or_ln896_54_fu_16485_p2 = (xor_ln896_137_fu_16479_p2 | xor_ln896_136_fu_16397_p2);

assign or_ln896_55_fu_14529_p2 = (xor_ln896_140_fu_14523_p2 | xor_ln896_139_fu_14431_p2);

assign or_ln896_56_fu_16677_p2 = (xor_ln896_142_fu_16671_p2 | xor_ln896_141_fu_16589_p2);

assign or_ln896_57_fu_14703_p2 = (xor_ln896_145_fu_14697_p2 | xor_ln896_144_fu_14605_p2);

assign or_ln896_58_fu_16851_p2 = (xor_ln896_147_fu_16845_p2 | xor_ln896_146_fu_16751_p2);

assign or_ln896_59_fu_18307_p2 = (xor_ln896_149_fu_18301_p2 | xor_ln896_148_fu_18207_p2);

assign or_ln896_5_fu_5454_p2 = (xor_ln896_11_fu_5448_p2 | xor_ln896_10_fu_5354_p2);

assign or_ln896_60_fu_14900_p2 = (xor_ln896_151_fu_14894_p2 | xor_ln896_150_fu_14802_p2);

assign or_ln896_61_fu_17088_p2 = (xor_ln896_153_fu_17082_p2 | xor_ln896_152_fu_16988_p2);

assign or_ln896_62_fu_18519_p2 = (xor_ln896_155_fu_18513_p2 | xor_ln896_154_fu_18419_p2);

assign or_ln896_6_fu_6144_p2 = (xor_ln896_13_fu_6138_p2 | xor_ln896_12_fu_6044_p2);

assign or_ln896_7_fu_6840_p2 = (xor_ln896_15_fu_6834_p2 | xor_ln896_14_fu_6740_p2);

assign or_ln896_8_fu_7552_p2 = (xor_ln896_17_fu_7546_p2 | xor_ln896_16_fu_7452_p2);

assign or_ln896_9_fu_8345_p2 = (xor_ln896_19_fu_8339_p2 | xor_ln896_18_fu_8245_p2);

assign or_ln896_fu_2123_p2 = (xor_ln896_fu_2025_p2 | xor_ln896_1_fu_2117_p2);

assign select_ln302_10_fu_2993_p3 = ((xor_ln302_10_fu_2979_p2[0:0] == 1'b1) ? select_ln346_27_fu_2985_p3 : add_ln813_10_fu_2953_p2);

assign select_ln302_11_fu_3063_p3 = ((xor_ln302_11_fu_3049_p2[0:0] == 1'b1) ? select_ln346_28_fu_3055_p3 : add_ln813_11_fu_3023_p2);

assign select_ln302_12_fu_3712_p3 = ((xor_ln302_12_fu_3698_p2[0:0] == 1'b1) ? select_ln346_29_fu_3704_p3 : add_ln813_12_fu_3672_p2);

assign select_ln302_13_fu_3782_p3 = ((xor_ln302_13_fu_3768_p2[0:0] == 1'b1) ? select_ln346_30_fu_3774_p3 : add_ln813_13_fu_3742_p2);

assign select_ln302_14_fu_4569_p3 = ((xor_ln302_14_fu_4555_p2[0:0] == 1'b1) ? select_ln346_31_fu_4561_p3 : add_ln813_14_fu_4529_p2);

assign select_ln302_15_fu_4639_p3 = ((xor_ln302_15_fu_4625_p2[0:0] == 1'b1) ? select_ln346_32_fu_4631_p3 : add_ln813_15_fu_4599_p2);

assign select_ln302_16_fu_5204_p3 = ((xor_ln302_16_fu_5190_p2[0:0] == 1'b1) ? select_ln346_33_fu_5196_p3 : add_ln813_16_fu_5164_p2);

assign select_ln302_17_fu_5274_p3 = ((xor_ln302_17_fu_5260_p2[0:0] == 1'b1) ? select_ln346_34_fu_5266_p3 : add_ln813_17_fu_5234_p2);

assign select_ln302_18_fu_1441_p3 = ((xor_ln302_18_fu_1427_p2[0:0] == 1'b1) ? select_ln346_18_fu_1433_p3 : add_ln813_1_fu_1401_p2);

assign select_ln302_19_fu_1589_p3 = ((xor_ln302_4_fu_1575_p2[0:0] == 1'b1) ? select_ln346_21_fu_1581_p3 : add_ln813_4_fu_1549_p2);

assign select_ln302_20_fu_1899_p3 = ((xor_ln302_6_fu_1885_p2[0:0] == 1'b1) ? select_ln346_23_fu_1891_p3 : add_ln813_6_fu_1859_p2);

assign select_ln302_21_fu_10332_p3 = ((xor_ln302_21_fu_10318_p2[0:0] == 1'b1) ? select_ln346_131_fu_10324_p3 : trunc_ln813_fu_10294_p1);

assign select_ln302_22_fu_9610_p3 = ((xor_ln302_22_fu_9596_p2[0:0] == 1'b1) ? select_ln346_132_fu_9602_p3 : trunc_ln813_18_fu_9572_p1);

assign select_ln302_23_fu_8709_p3 = ((xor_ln302_23_fu_8695_p2[0:0] == 1'b1) ? select_ln346_133_fu_8701_p3 : trunc_ln813_19_fu_8671_p1);

assign select_ln302_24_fu_18621_p3 = ((xor_ln302_24_fu_18607_p2[0:0] == 1'b1) ? select_ln346_248_fu_18613_p3 : add_ln813_18_fu_18581_p2);

assign select_ln302_25_fu_18692_p3 = ((xor_ln302_25_fu_18678_p2[0:0] == 1'b1) ? select_ln346_249_fu_18684_p3 : add_ln813_19_fu_18652_p2);

assign select_ln302_26_fu_18797_p3 = ((xor_ln302_26_fu_18783_p2[0:0] == 1'b1) ? select_ln346_250_fu_18789_p3 : add_ln813_20_fu_18757_p2);

assign select_ln302_27_fu_18868_p3 = ((xor_ln302_27_fu_18854_p2[0:0] == 1'b1) ? select_ln346_251_fu_18860_p3 : add_ln813_21_fu_18828_p2);

assign select_ln302_28_fu_18973_p3 = ((xor_ln302_28_fu_18959_p2[0:0] == 1'b1) ? select_ln346_252_fu_18965_p3 : add_ln813_22_fu_18933_p2);

assign select_ln302_29_fu_19044_p3 = ((xor_ln302_29_fu_19030_p2[0:0] == 1'b1) ? select_ln346_253_fu_19036_p3 : add_ln813_23_fu_19004_p2);

assign select_ln302_2_fu_1519_p3 = ((xor_ln302_19_fu_1505_p2[0:0] == 1'b1) ? select_ln346_19_fu_1511_p3 : add_ln813_2_fu_1479_p2);

assign select_ln302_30_fu_19149_p3 = ((xor_ln302_30_fu_19135_p2[0:0] == 1'b1) ? select_ln346_254_fu_19141_p3 : add_ln813_24_fu_19109_p2);

assign select_ln302_31_fu_19220_p3 = ((xor_ln302_31_fu_19206_p2[0:0] == 1'b1) ? select_ln346_255_fu_19212_p3 : add_ln813_25_fu_19180_p2);

assign select_ln302_32_fu_19325_p3 = ((xor_ln302_32_fu_19311_p2[0:0] == 1'b1) ? select_ln346_256_fu_19317_p3 : add_ln813_26_fu_19285_p2);

assign select_ln302_33_fu_19396_p3 = ((xor_ln302_33_fu_19382_p2[0:0] == 1'b1) ? select_ln346_257_fu_19388_p3 : add_ln813_27_fu_19356_p2);

assign select_ln302_34_fu_19501_p3 = ((xor_ln302_34_fu_19487_p2[0:0] == 1'b1) ? select_ln346_258_fu_19493_p3 : add_ln813_28_fu_19461_p2);

assign select_ln302_35_fu_19572_p3 = ((xor_ln302_35_fu_19558_p2[0:0] == 1'b1) ? select_ln346_259_fu_19564_p3 : add_ln813_29_fu_19532_p2);

assign select_ln302_36_fu_19677_p3 = ((xor_ln302_36_fu_19663_p2[0:0] == 1'b1) ? select_ln346_260_fu_19669_p3 : add_ln813_30_fu_19637_p2);

assign select_ln302_37_fu_19748_p3 = ((xor_ln302_37_fu_19734_p2[0:0] == 1'b1) ? select_ln346_261_fu_19740_p3 : add_ln813_31_fu_19708_p2);

assign select_ln302_38_fu_19853_p3 = ((xor_ln302_38_fu_19839_p2[0:0] == 1'b1) ? select_ln346_262_fu_19845_p3 : add_ln813_32_fu_19813_p2);

assign select_ln302_39_fu_19924_p3 = ((xor_ln302_39_fu_19910_p2[0:0] == 1'b1) ? select_ln346_263_fu_19916_p3 : add_ln813_33_fu_19884_p2);

assign select_ln302_3_fu_1671_p3 = ((xor_ln302_20_fu_1657_p2[0:0] == 1'b1) ? select_ln346_20_fu_1663_p3 : add_ln813_3_fu_1631_p2);

assign select_ln302_40_fu_20029_p3 = ((xor_ln302_40_fu_20015_p2[0:0] == 1'b1) ? select_ln346_264_fu_20021_p3 : add_ln813_34_fu_19989_p2);

assign select_ln302_41_fu_20100_p3 = ((xor_ln302_41_fu_20086_p2[0:0] == 1'b1) ? select_ln346_265_fu_20092_p3 : add_ln813_35_fu_20060_p2);

assign select_ln302_42_fu_20203_p3 = ((xor_ln302_42_fu_20189_p2[0:0] == 1'b1) ? select_ln346_266_fu_20195_p3 : add_ln813_36_fu_20164_p2);

assign select_ln302_43_fu_20272_p3 = ((xor_ln302_43_fu_20258_p2[0:0] == 1'b1) ? select_ln346_267_fu_20264_p3 : add_ln813_37_fu_20233_p2);

assign select_ln302_44_fu_20341_p3 = ((xor_ln302_44_fu_20327_p2[0:0] == 1'b1) ? select_ln346_268_fu_20333_p3 : add_ln813_38_fu_20302_p2);

assign select_ln302_45_fu_20410_p3 = ((xor_ln302_45_fu_20396_p2[0:0] == 1'b1) ? select_ln346_269_fu_20402_p3 : add_ln813_39_fu_20371_p2);

assign select_ln302_46_fu_20479_p3 = ((xor_ln302_46_fu_20465_p2[0:0] == 1'b1) ? select_ln346_270_fu_20471_p3 : add_ln813_40_fu_20440_p2);

assign select_ln302_47_fu_20548_p3 = ((xor_ln302_47_fu_20534_p2[0:0] == 1'b1) ? select_ln346_271_fu_20540_p3 : add_ln813_41_fu_20509_p2);

assign select_ln302_48_fu_20617_p3 = ((xor_ln302_48_fu_20603_p2[0:0] == 1'b1) ? select_ln346_272_fu_20609_p3 : add_ln813_42_fu_20578_p2);

assign select_ln302_49_fu_20686_p3 = ((xor_ln302_49_fu_20672_p2[0:0] == 1'b1) ? select_ln346_273_fu_20678_p3 : add_ln813_43_fu_20647_p2);

assign select_ln302_50_fu_20755_p3 = ((xor_ln302_50_fu_20741_p2[0:0] == 1'b1) ? select_ln346_274_fu_20747_p3 : add_ln813_44_fu_20716_p2);

assign select_ln302_51_fu_20824_p3 = ((xor_ln302_51_fu_20810_p2[0:0] == 1'b1) ? select_ln346_275_fu_20816_p3 : add_ln813_45_fu_20785_p2);

assign select_ln302_52_fu_20893_p3 = ((xor_ln302_52_fu_20879_p2[0:0] == 1'b1) ? select_ln346_276_fu_20885_p3 : add_ln813_46_fu_20854_p2);

assign select_ln302_53_fu_20962_p3 = ((xor_ln302_53_fu_20948_p2[0:0] == 1'b1) ? select_ln346_277_fu_20954_p3 : add_ln813_47_fu_20923_p2);

assign select_ln302_54_fu_21031_p3 = ((xor_ln302_54_fu_21017_p2[0:0] == 1'b1) ? select_ln346_278_fu_21023_p3 : add_ln813_48_fu_20992_p2);

assign select_ln302_55_fu_21100_p3 = ((xor_ln302_55_fu_21086_p2[0:0] == 1'b1) ? select_ln346_279_fu_21092_p3 : add_ln813_49_fu_21061_p2);

assign select_ln302_56_fu_21169_p3 = ((xor_ln302_56_fu_21155_p2[0:0] == 1'b1) ? select_ln346_280_fu_21161_p3 : add_ln813_50_fu_21130_p2);

assign select_ln302_57_fu_21238_p3 = ((xor_ln302_57_fu_21224_p2[0:0] == 1'b1) ? select_ln346_281_fu_21230_p3 : add_ln813_51_fu_21199_p2);

assign select_ln302_58_fu_21307_p3 = ((xor_ln302_58_fu_21293_p2[0:0] == 1'b1) ? select_ln346_282_fu_21299_p3 : add_ln813_52_fu_21268_p2);

assign select_ln302_59_fu_21376_p3 = ((xor_ln302_59_fu_21362_p2[0:0] == 1'b1) ? select_ln346_283_fu_21368_p3 : add_ln813_53_fu_21337_p2);

assign select_ln302_5_fu_1741_p3 = ((xor_ln302_5_fu_1727_p2[0:0] == 1'b1) ? select_ln346_22_fu_1733_p3 : add_ln813_5_fu_1701_p2);

assign select_ln302_7_fu_1969_p3 = ((xor_ln302_7_fu_1955_p2[0:0] == 1'b1) ? select_ln346_24_fu_1961_p3 : add_ln813_7_fu_1929_p2);

assign select_ln302_8_fu_2240_p3 = ((xor_ln302_8_fu_2226_p2[0:0] == 1'b1) ? select_ln346_25_fu_2232_p3 : add_ln813_8_fu_2200_p2);

assign select_ln302_9_fu_2310_p3 = ((xor_ln302_9_fu_2296_p2[0:0] == 1'b1) ? select_ln346_26_fu_2302_p3 : add_ln813_9_fu_2270_p2);

assign select_ln302_fu_1371_p3 = ((xor_ln302_fu_1357_p2[0:0] == 1'b1) ? select_ln346_fu_1363_p3 : add_ln813_fu_1331_p2);

assign select_ln346_100_fu_9499_p3 = ((or_ln346_23_reg_23135[0:0] == 1'b1) ? select_ln346_99_fu_9492_p3 : add_ln377_23_reg_23125);

assign select_ln346_101_fu_9533_p3 = ((and_ln895_68_fu_9527_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_102_fu_9547_p3 = ((xor_ln346_9_fu_9541_p2[0:0] == 1'b1) ? select_ln346_101_fu_9533_p3 : select_ln346_100_fu_9499_p3);

assign select_ln346_103_fu_2915_p3 = ((and_ln895_69_fu_2879_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_104_fu_2923_p3 = ((or_ln346_24_fu_2909_p2[0:0] == 1'b1) ? select_ln346_103_fu_2915_p3 : add_ln377_24_fu_2779_p2);

assign select_ln346_105_fu_4288_p3 = ((and_ln895_70_reg_22620[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_106_fu_4300_p3 = ((or_ln346_25_fu_4295_p2[0:0] == 1'b1) ? select_ln346_105_fu_4288_p3 : add_ln377_25_reg_22605);

assign select_ln346_107_fu_4335_p3 = ((and_ln895_71_fu_4329_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_108_fu_4349_p3 = ((xor_ln346_10_fu_4343_p2[0:0] == 1'b1) ? select_ln346_107_fu_4335_p3 : select_ln346_106_fu_4300_p3);

assign select_ln346_109_fu_4385_p3 = ((and_ln895_72_fu_4379_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_110_fu_4399_p3 = ((xor_ln346_11_fu_4393_p2[0:0] == 1'b1) ? select_ln346_109_fu_4385_p3 : select_ln346_108_fu_4349_p3);

assign select_ln346_111_fu_4435_p3 = ((and_ln895_73_fu_4429_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_112_fu_4449_p3 = ((xor_ln346_12_fu_4443_p2[0:0] == 1'b1) ? select_ln346_111_fu_4435_p3 : select_ln346_110_fu_4399_p3);

assign select_ln346_113_fu_4491_p3 = ((and_ln895_74_fu_4479_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_114_fu_4499_p3 = ((xor_ln346_13_fu_4485_p2[0:0] == 1'b1) ? select_ln346_113_fu_4491_p3 : select_ln346_112_fu_4449_p3);

assign select_ln346_115_fu_6457_p3 = ((and_ln895_75_reg_22865[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_116_fu_6464_p3 = ((or_ln346_26_fu_6452_p2[0:0] == 1'b1) ? select_ln346_115_fu_6457_p3 : add_ln377_26_reg_22850);

assign select_ln346_117_fu_7109_p3 = ((and_ln895_76_reg_22937[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_118_fu_7116_p3 = ((or_ln346_27_reg_22942[0:0] == 1'b1) ? select_ln346_117_fu_7109_p3 : add_ln377_27_reg_22932);

assign select_ln346_119_fu_7150_p3 = ((and_ln895_77_fu_7144_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_120_fu_7164_p3 = ((xor_ln346_14_fu_7158_p2[0:0] == 1'b1) ? select_ln346_119_fu_7150_p3 : select_ln346_118_fu_7116_p3);

assign select_ln346_121_fu_7206_p3 = ((and_ln895_78_fu_7194_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_122_fu_7214_p3 = ((xor_ln346_15_fu_7200_p2[0:0] == 1'b1) ? select_ln346_121_fu_7206_p3 : select_ln346_120_fu_7164_p3);

assign select_ln346_123_fu_7853_p3 = ((and_ln895_79_reg_22992[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_124_fu_7865_p3 = ((or_ln346_28_fu_7860_p2[0:0] == 1'b1) ? select_ln346_123_fu_7853_p3 : add_ln377_28_reg_22977);

assign select_ln346_125_fu_7900_p3 = ((and_ln895_80_fu_7894_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_126_fu_7914_p3 = ((xor_ln346_16_fu_7908_p2[0:0] == 1'b1) ? select_ln346_125_fu_7900_p3 : select_ln346_124_fu_7865_p3);

assign select_ln346_127_fu_7956_p3 = ((and_ln895_81_fu_7944_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_128_fu_7964_p3 = ((xor_ln346_17_fu_7950_p2[0:0] == 1'b1) ? select_ln346_127_fu_7956_p3 : select_ln346_126_fu_7914_p3);

assign select_ln346_129_fu_8635_p3 = ((and_ln895_82_reg_23058[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_130_fu_8647_p3 = ((or_ln346_29_fu_8642_p2[0:0] == 1'b1) ? select_ln346_129_fu_8635_p3 : add_ln377_29_reg_23043);

assign select_ln346_131_fu_10324_p3 = ((and_ln895_83_fu_10312_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_132_fu_9602_p3 = ((and_ln895_84_fu_9590_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_133_fu_8701_p3 = ((and_ln895_85_fu_8689_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_134_fu_10540_p3 = ((and_ln895_86_fu_10504_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_135_fu_10548_p3 = ((or_ln346_30_fu_10534_p2[0:0] == 1'b1) ? select_ln346_134_fu_10540_p3 : add_ln377_30_fu_10404_p2);

assign select_ln346_136_fu_11103_p3 = ((and_ln895_87_fu_11067_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_137_fu_11111_p3 = ((or_ln346_31_fu_11097_p2[0:0] == 1'b1) ? select_ln346_136_fu_11103_p3 : add_ln377_31_fu_10965_p2);

assign select_ln346_138_fu_12180_p3 = ((and_ln895_88_reg_23330[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_139_fu_12187_p3 = ((or_ln346_32_reg_23335[0:0] == 1'b1) ? select_ln346_138_fu_12180_p3 : add_ln377_32_reg_23325);

assign select_ln346_140_fu_11122_p3 = ((and_ln895_89_reg_23275[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_141_fu_11129_p3 = ((or_ln346_33_reg_23280[0:0] == 1'b1) ? select_ln346_140_fu_11122_p3 : sext_ln856_fu_11119_p1);

assign select_ln346_142_fu_11333_p3 = ((and_ln895_90_fu_11297_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_143_fu_11341_p3 = ((or_ln346_34_fu_11327_p2[0:0] == 1'b1) ? select_ln346_142_fu_11333_p3 : add_ln377_34_fu_11195_p2);

assign select_ln346_144_fu_12199_p3 = ((and_ln895_91_reg_23345[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_145_fu_12206_p3 = ((or_ln346_35_reg_23350[0:0] == 1'b1) ? select_ln346_144_fu_12199_p3 : add_ln377_35_reg_23340);

assign select_ln346_146_fu_11369_p3 = ((and_ln895_92_reg_23290[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_147_fu_11376_p3 = ((or_ln346_36_reg_23295[0:0] == 1'b1) ? select_ln346_146_fu_11369_p3 : sext_ln856_1_fu_11349_p1);

assign select_ln346_148_fu_11974_p3 = ((and_ln895_93_reg_23315[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_149_fu_11981_p3 = ((or_ln346_37_reg_23320[0:0] == 1'b1) ? select_ln346_148_fu_11974_p3 : add_ln377_37_reg_23310);

assign select_ln346_150_fu_12524_p3 = ((and_ln895_94_reg_23360[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_151_fu_12531_p3 = ((or_ln346_38_reg_23365[0:0] == 1'b1) ? select_ln346_150_fu_12524_p3 : add_ln377_38_reg_23355);

assign select_ln346_152_fu_14931_p3 = ((and_ln895_95_reg_23455[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_153_fu_14938_p3 = ((or_ln346_39_reg_23460[0:0] == 1'b1) ? select_ln346_152_fu_14931_p3 : add_ln377_39_reg_23450);

assign select_ln346_154_fu_14972_p3 = ((and_ln895_96_fu_14966_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_155_fu_14986_p3 = ((xor_ln346_18_fu_14980_p2[0:0] == 1'b1) ? select_ln346_154_fu_14972_p3 : select_ln346_153_fu_14938_p3);

assign select_ln346_156_fu_15022_p3 = ((and_ln895_97_fu_15016_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_157_fu_15036_p3 = ((xor_ln346_19_fu_15030_p2[0:0] == 1'b1) ? select_ln346_156_fu_15022_p3 : select_ln346_155_fu_14986_p3);

assign select_ln346_158_fu_15048_p3 = ((and_ln895_98_reg_23470[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_159_fu_15055_p3 = ((or_ln346_40_reg_23475[0:0] == 1'b1) ? select_ln346_158_fu_15048_p3 : sext_ln856_2_fu_15045_p1);

assign select_ln346_160_fu_15090_p3 = ((and_ln895_99_fu_15084_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_161_fu_15104_p3 = ((xor_ln346_20_fu_15098_p2[0:0] == 1'b1) ? select_ln346_160_fu_15090_p3 : select_ln346_159_fu_15055_p3);

assign select_ln346_162_fu_15140_p3 = ((and_ln895_100_fu_15134_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_163_fu_15154_p3 = ((xor_ln346_21_fu_15148_p2[0:0] == 1'b1) ? select_ln346_162_fu_15140_p3 : select_ln346_161_fu_15104_p3);

assign select_ln346_164_fu_13625_p3 = ((and_ln895_101_fu_13589_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_165_fu_13633_p3 = ((or_ln346_41_fu_13619_p2[0:0] == 1'b1) ? select_ln346_164_fu_13625_p3 : add_ln377_41_fu_13489_p2);

assign select_ln346_166_fu_17154_p3 = ((and_ln895_102_reg_23629[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_167_fu_17166_p3 = ((or_ln346_42_fu_17161_p2[0:0] == 1'b1) ? select_ln346_166_fu_17154_p3 : add_ln377_42_reg_23614);

assign select_ln346_168_fu_17201_p3 = ((and_ln895_103_fu_17195_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_169_fu_17215_p3 = ((xor_ln346_22_fu_17209_p2[0:0] == 1'b1) ? select_ln346_168_fu_17201_p3 : select_ln346_167_fu_17166_p3);

assign select_ln346_170_fu_15336_p3 = ((and_ln895_104_reg_23490[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_171_fu_15343_p3 = ((or_ln346_43_reg_23495[0:0] == 1'b1) ? select_ln346_170_fu_15336_p3 : sext_ln856_3_fu_15333_p1);

assign select_ln346_172_fu_17242_p3 = ((and_ln895_105_reg_23665[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_173_fu_17254_p3 = ((or_ln346_44_fu_17249_p2[0:0] == 1'b1) ? select_ln346_172_fu_17242_p3 : add_ln377_44_reg_23650);

assign select_ln346_174_fu_17289_p3 = ((and_ln895_106_fu_17283_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_175_fu_17303_p3 = ((xor_ln346_23_fu_17297_p2[0:0] == 1'b1) ? select_ln346_174_fu_17289_p3 : select_ln346_173_fu_17254_p3);

assign select_ln346_176_fu_13989_p3 = ((and_ln895_107_fu_13953_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_177_fu_13997_p3 = ((or_ln346_45_fu_13983_p2[0:0] == 1'b1) ? select_ln346_176_fu_13989_p3 : add_ln377_45_fu_13853_p2);

assign select_ln346_178_fu_15717_p3 = ((and_ln895_108_fu_15681_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_179_fu_15725_p3 = ((or_ln346_46_fu_15711_p2[0:0] == 1'b1) ? select_ln346_178_fu_15717_p3 : add_ln377_46_fu_15579_p2);

assign select_ln346_180_fu_17497_p3 = ((and_ln895_109_fu_17467_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_181_fu_17511_p3 = ((or_ln346_47_fu_17505_p2[0:0] == 1'b1) ? select_ln346_180_fu_17497_p3 : add_ln377_47_fu_17365_p2);

assign select_ln346_182_fu_15743_p3 = ((and_ln895_110_reg_23521[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_183_fu_15750_p3 = ((or_ln346_48_reg_23526[0:0] == 1'b1) ? select_ln346_182_fu_15743_p3 : sext_ln856_4_fu_15740_p1);

assign select_ln346_184_fu_15954_p3 = ((and_ln895_111_fu_15918_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_185_fu_15962_p3 = ((or_ln346_49_fu_15948_p2[0:0] == 1'b1) ? select_ln346_184_fu_15954_p3 : add_ln377_49_fu_15816_p2);

assign select_ln346_186_fu_17709_p3 = ((and_ln895_112_fu_17679_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_187_fu_17723_p3 = ((or_ln346_50_fu_17717_p2[0:0] == 1'b1) ? select_ln346_186_fu_17709_p3 : add_ln377_50_fu_17577_p2);

assign select_ln346_188_fu_17731_p3 = ((and_ln895_113_reg_23713[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_189_fu_17738_p3 = ((or_ln346_51_reg_23718[0:0] == 1'b1) ? select_ln346_188_fu_17731_p3 : add_ln377_51_reg_23708);

assign select_ln346_18_fu_1433_p3 = ((and_ln895_18_fu_1421_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_190_fu_17772_p3 = ((and_ln895_114_fu_17766_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_191_fu_17786_p3 = ((xor_ln346_24_fu_17780_p2[0:0] == 1'b1) ? select_ln346_190_fu_17772_p3 : select_ln346_189_fu_17738_p3);

assign select_ln346_192_fu_17822_p3 = ((and_ln895_115_fu_17816_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_193_fu_17836_p3 = ((xor_ln346_25_fu_17830_p2[0:0] == 1'b1) ? select_ln346_192_fu_17822_p3 : select_ln346_191_fu_17786_p3);

assign select_ln346_194_fu_17848_p3 = ((and_ln895_116_reg_23728[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_195_fu_17855_p3 = ((or_ln346_52_reg_23733[0:0] == 1'b1) ? select_ln346_194_fu_17848_p3 : sext_ln856_5_fu_17845_p1);

assign select_ln346_196_fu_17890_p3 = ((and_ln895_117_fu_17884_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_197_fu_17904_p3 = ((xor_ln346_26_fu_17898_p2[0:0] == 1'b1) ? select_ln346_196_fu_17890_p3 : select_ln346_195_fu_17855_p3);

assign select_ln346_198_fu_17940_p3 = ((and_ln895_118_fu_17934_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_199_fu_17954_p3 = ((xor_ln346_27_fu_17948_p2[0:0] == 1'b1) ? select_ln346_198_fu_17940_p3 : select_ln346_197_fu_17904_p3);

assign select_ln346_19_fu_1511_p3 = ((and_ln895_19_fu_1499_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_200_fu_14363_p3 = ((and_ln895_119_fu_14327_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_201_fu_14371_p3 = ((or_ln346_53_fu_14357_p2[0:0] == 1'b1) ? select_ln346_200_fu_14363_p3 : add_ln377_53_fu_14227_p2);

assign select_ln346_202_fu_17982_p3 = ((and_ln895_120_reg_23763[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_203_fu_17994_p3 = ((or_ln346_54_fu_17989_p2[0:0] == 1'b1) ? select_ln346_202_fu_17982_p3 : add_ln377_54_reg_23748);

assign select_ln346_204_fu_18029_p3 = ((and_ln895_121_fu_18023_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_205_fu_18043_p3 = ((xor_ln346_28_fu_18037_p2[0:0] == 1'b1) ? select_ln346_204_fu_18029_p3 : select_ln346_203_fu_17994_p3);

assign select_ln346_206_fu_16494_p3 = ((and_ln895_122_reg_23552[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_207_fu_16501_p3 = ((or_ln346_55_reg_23557[0:0] == 1'b1) ? select_ln346_206_fu_16494_p3 : sext_ln856_6_fu_16491_p1);

assign select_ln346_208_fu_18070_p3 = ((and_ln895_123_reg_23799[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_209_fu_18082_p3 = ((or_ln346_56_fu_18077_p2[0:0] == 1'b1) ? select_ln346_208_fu_18070_p3 : add_ln377_56_reg_23784);

assign select_ln346_20_fu_1663_p3 = ((and_ln895_20_fu_1651_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_210_fu_18117_p3 = ((and_ln895_124_fu_18111_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_211_fu_18131_p3 = ((xor_ln346_29_fu_18125_p2[0:0] == 1'b1) ? select_ln346_210_fu_18117_p3 : select_ln346_209_fu_18082_p3);

assign select_ln346_212_fu_14727_p3 = ((and_ln895_125_fu_14691_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_213_fu_14735_p3 = ((or_ln346_57_fu_14721_p2[0:0] == 1'b1) ? select_ln346_212_fu_14727_p3 : add_ln377_57_fu_14591_p2);

assign select_ln346_214_fu_16875_p3 = ((and_ln895_126_fu_16839_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_215_fu_16883_p3 = ((or_ln346_58_fu_16869_p2[0:0] == 1'b1) ? select_ln346_214_fu_16875_p3 : add_ln377_58_fu_16737_p2);

assign select_ln346_216_fu_18325_p3 = ((and_ln895_127_fu_18295_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_217_fu_18339_p3 = ((or_ln346_59_fu_18333_p2[0:0] == 1'b1) ? select_ln346_216_fu_18325_p3 : add_ln377_59_fu_18193_p2);

assign select_ln346_218_fu_16901_p3 = ((and_ln895_128_reg_23583[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_219_fu_16908_p3 = ((or_ln346_60_reg_23588[0:0] == 1'b1) ? select_ln346_218_fu_16901_p3 : sext_ln856_7_fu_16898_p1);

assign select_ln346_21_fu_1581_p3 = ((and_ln895_21_fu_1569_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_220_fu_17112_p3 = ((and_ln895_129_fu_17076_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_221_fu_17120_p3 = ((or_ln346_61_fu_17106_p2[0:0] == 1'b1) ? select_ln346_220_fu_17112_p3 : add_ln377_61_fu_16974_p2);

assign select_ln346_222_fu_18537_p3 = ((and_ln895_130_fu_18507_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_223_fu_18551_p3 = ((or_ln346_62_fu_18545_p2[0:0] == 1'b1) ? select_ln346_222_fu_18537_p3 : add_ln377_62_fu_18405_p2);

assign select_ln346_224_fu_12268_p3 = ((and_ln895_131_fu_12262_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_225_fu_12282_p3 = ((xor_ln346_30_fu_12276_p2[0:0] == 1'b1) ? select_ln346_224_fu_12268_p3 : select_ln346_139_fu_12187_p3);

assign select_ln346_226_fu_12318_p3 = ((and_ln895_132_fu_12312_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_227_fu_12332_p3 = ((xor_ln346_31_fu_12326_p2[0:0] == 1'b1) ? select_ln346_226_fu_12318_p3 : select_ln346_225_fu_12282_p3);

assign select_ln346_228_fu_12368_p3 = ((and_ln895_133_fu_12362_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_229_fu_12382_p3 = ((xor_ln346_32_fu_12376_p2[0:0] == 1'b1) ? select_ln346_228_fu_12368_p3 : select_ln346_227_fu_12332_p3);

assign select_ln346_22_fu_1733_p3 = ((and_ln895_22_fu_1721_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_230_fu_12451_p3 = ((and_ln895_134_fu_12427_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_231_fu_12465_p3 = ((or_ln346_63_fu_12459_p2[0:0] == 1'b1) ? select_ln346_230_fu_12451_p3 : select_ln346_145_fu_12206_p3);

assign select_ln346_232_fu_12501_p3 = ((and_ln895_135_fu_12495_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_233_fu_12515_p3 = ((xor_ln346_33_fu_12509_p2[0:0] == 1'b1) ? select_ln346_232_fu_12501_p3 : select_ln346_231_fu_12465_p3);

assign select_ln346_234_fu_12608_p3 = ((and_ln895_136_fu_12584_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_235_fu_12622_p3 = ((or_ln346_64_fu_12616_p2[0:0] == 1'b1) ? select_ln346_234_fu_12608_p3 : select_ln346_151_fu_12531_p3);

assign select_ln346_236_fu_12718_p3 = ((and_ln895_137_fu_12694_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_237_fu_12732_p3 = ((or_ln346_65_fu_12726_p2[0:0] == 1'b1) ? select_ln346_236_fu_12718_p3 : trunc_ln818_62_fu_12656_p4);

assign select_ln346_238_fu_12768_p3 = ((and_ln895_138_fu_12762_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_239_fu_12782_p3 = ((xor_ln346_34_fu_12776_p2[0:0] == 1'b1) ? select_ln346_238_fu_12768_p3 : select_ln346_237_fu_12732_p3);

assign select_ln346_23_fu_1891_p3 = ((and_ln895_23_fu_1879_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_240_fu_12818_p3 = ((and_ln895_139_fu_12812_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_241_fu_12832_p3 = ((xor_ln346_35_fu_12826_p2[0:0] == 1'b1) ? select_ln346_240_fu_12818_p3 : select_ln346_239_fu_12782_p3);

assign select_ln346_242_fu_12939_p3 = ((and_ln895_140_fu_12915_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_243_fu_12953_p3 = ((or_ln346_66_fu_12947_p2[0:0] == 1'b1) ? select_ln346_242_fu_12939_p3 : trunc_ln818_63_fu_12877_p4);

assign select_ln346_244_fu_12989_p3 = ((and_ln895_141_fu_12983_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_245_fu_13003_p3 = ((xor_ln346_36_fu_12997_p2[0:0] == 1'b1) ? select_ln346_244_fu_12989_p3 : select_ln346_243_fu_12953_p3);

assign select_ln346_246_fu_13088_p3 = ((and_ln895_142_fu_13064_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_247_fu_13102_p3 = ((or_ln346_67_fu_13096_p2[0:0] == 1'b1) ? select_ln346_246_fu_13088_p3 : trunc_ln818_64_fu_13026_p4);

assign select_ln346_248_fu_18613_p3 = ((and_ln895_143_fu_18601_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_249_fu_18684_p3 = ((and_ln895_144_fu_18672_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_24_fu_1961_p3 = ((and_ln895_24_fu_1949_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_250_fu_18789_p3 = ((and_ln895_145_fu_18777_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_251_fu_18860_p3 = ((and_ln895_146_fu_18848_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_252_fu_18965_p3 = ((and_ln895_147_fu_18953_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_253_fu_19036_p3 = ((and_ln895_148_fu_19024_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_254_fu_19141_p3 = ((and_ln895_149_fu_19129_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_255_fu_19212_p3 = ((and_ln895_150_fu_19200_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_256_fu_19317_p3 = ((and_ln895_151_fu_19305_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_257_fu_19388_p3 = ((and_ln895_152_fu_19376_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_258_fu_19493_p3 = ((and_ln895_153_fu_19481_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_259_fu_19564_p3 = ((and_ln895_154_fu_19552_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_25_fu_2232_p3 = ((and_ln895_25_fu_2220_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_260_fu_19669_p3 = ((and_ln895_155_fu_19657_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_261_fu_19740_p3 = ((and_ln895_156_fu_19728_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_262_fu_19845_p3 = ((and_ln895_157_fu_19833_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_263_fu_19916_p3 = ((and_ln895_158_fu_19904_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_264_fu_20021_p3 = ((and_ln895_159_fu_20009_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_265_fu_20092_p3 = ((and_ln895_160_fu_20080_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_266_fu_20195_p3 = ((and_ln895_161_fu_20183_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_267_fu_20264_p3 = ((and_ln895_162_fu_20252_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_268_fu_20333_p3 = ((and_ln895_163_fu_20321_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_269_fu_20402_p3 = ((and_ln895_164_fu_20390_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_26_fu_2302_p3 = ((and_ln895_26_fu_2290_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_270_fu_20471_p3 = ((and_ln895_165_fu_20459_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_271_fu_20540_p3 = ((and_ln895_166_fu_20528_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_272_fu_20609_p3 = ((and_ln895_167_fu_20597_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_273_fu_20678_p3 = ((and_ln895_168_fu_20666_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_274_fu_20747_p3 = ((and_ln895_169_fu_20735_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_275_fu_20816_p3 = ((and_ln895_170_fu_20804_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_276_fu_20885_p3 = ((and_ln895_171_fu_20873_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_277_fu_20954_p3 = ((and_ln895_172_fu_20942_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_278_fu_21023_p3 = ((and_ln895_173_fu_21011_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_279_fu_21092_p3 = ((and_ln895_174_fu_21080_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_27_fu_2985_p3 = ((and_ln895_27_fu_2973_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_280_fu_21161_p3 = ((and_ln895_175_fu_21149_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_281_fu_21230_p3 = ((and_ln895_176_fu_21218_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_282_fu_21299_p3 = ((and_ln895_177_fu_21287_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_283_fu_21368_p3 = ((and_ln895_178_fu_21356_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_28_fu_3055_p3 = ((and_ln895_28_fu_3043_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_29_fu_3704_p3 = ((and_ln895_29_fu_3692_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_30_fu_3774_p3 = ((and_ln895_30_fu_3762_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_31_fu_4561_p3 = ((and_ln895_31_fu_4549_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_32_fu_4631_p3 = ((and_ln895_32_fu_4619_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_33_fu_5196_p3 = ((and_ln895_33_fu_5184_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_34_fu_5266_p3 = ((and_ln895_34_fu_5254_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_35_fu_2147_p3 = ((and_ln895_35_fu_2111_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_36_fu_2155_p3 = ((or_ln346_fu_2141_p2[0:0] == 1'b1) ? select_ln346_35_fu_2147_p3 : add_ln377_fu_2011_p2);

assign select_ln346_37_fu_2514_p3 = ((and_ln895_36_fu_2478_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_38_fu_2522_p3 = ((or_ln346_1_fu_2508_p2[0:0] == 1'b1) ? select_ln346_37_fu_2514_p3 : add_ln377_1_fu_2376_p2);

assign select_ln346_39_fu_3263_p3 = ((and_ln895_37_fu_3227_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_40_fu_3271_p3 = ((or_ln346_2_fu_3257_p2[0:0] == 1'b1) ? select_ln346_39_fu_3263_p3 : add_ln377_2_fu_3125_p2);

assign select_ln346_41_fu_4647_p3 = ((and_ln895_38_reg_22636[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_42_fu_4654_p3 = ((or_ln346_3_reg_22641[0:0] == 1'b1) ? select_ln346_41_fu_4647_p3 : add_ln377_3_reg_22631);

assign select_ln346_43_fu_4857_p3 = ((and_ln895_39_fu_4821_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_44_fu_4865_p3 = ((or_ln346_4_fu_4851_p2[0:0] == 1'b1) ? select_ln346_43_fu_4857_p3 : add_ln377_4_fu_4719_p2);

assign select_ln346_45_fu_5478_p3 = ((and_ln895_40_fu_5442_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_46_fu_5486_p3 = ((or_ln346_5_fu_5472_p2[0:0] == 1'b1) ? select_ln346_45_fu_5478_p3 : add_ln377_5_fu_5340_p2);

assign select_ln346_47_fu_6168_p3 = ((and_ln895_41_fu_6132_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_48_fu_6176_p3 = ((or_ln346_6_fu_6162_p2[0:0] == 1'b1) ? select_ln346_47_fu_6168_p3 : add_ln377_6_fu_6030_p2);

assign select_ln346_49_fu_6864_p3 = ((and_ln895_42_fu_6828_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_50_fu_6872_p3 = ((or_ln346_7_fu_6858_p2[0:0] == 1'b1) ? select_ln346_49_fu_6864_p3 : add_ln377_7_fu_6726_p2);

assign select_ln346_51_fu_7576_p3 = ((and_ln895_43_fu_7540_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_52_fu_7584_p3 = ((or_ln346_8_fu_7570_p2[0:0] == 1'b1) ? select_ln346_51_fu_7576_p3 : add_ln377_8_fu_7438_p2);

assign select_ln346_53_fu_8773_p3 = ((and_ln895_44_reg_23074[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_54_fu_8780_p3 = ((or_ln346_9_reg_23079[0:0] == 1'b1) ? select_ln346_53_fu_8773_p3 : add_ln377_9_reg_23069);

assign select_ln346_55_fu_8983_p3 = ((and_ln895_45_fu_8947_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_56_fu_8991_p3 = ((or_ln346_10_fu_8977_p2[0:0] == 1'b1) ? select_ln346_55_fu_8983_p3 : add_ln377_10_fu_8845_p2);

assign select_ln346_57_fu_9656_p3 = ((and_ln895_46_reg_23145[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_58_fu_9663_p3 = ((or_ln346_11_reg_23150[0:0] == 1'b1) ? select_ln346_57_fu_9656_p3 : add_ln377_11_reg_23140);

assign select_ln346_59_fu_9867_p3 = ((and_ln895_47_reg_23181[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_60_fu_9874_p3 = ((or_ln346_12_reg_23186[0:0] == 1'b1) ? select_ln346_59_fu_9867_p3 : add_ln377_12_reg_23176);

assign select_ln346_61_fu_9908_p3 = ((and_ln895_48_fu_9902_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_62_fu_9922_p3 = ((xor_ln346_fu_9916_p2[0:0] == 1'b1) ? select_ln346_61_fu_9908_p3 : select_ln346_60_fu_9874_p3);

assign select_ln346_63_fu_9964_p3 = ((and_ln895_49_fu_9952_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_64_fu_9972_p3 = ((xor_ln346_1_fu_9958_p2[0:0] == 1'b1) ? select_ln346_63_fu_9964_p3 : select_ln346_62_fu_9922_p3);

assign select_ln346_65_fu_10164_p3 = ((and_ln895_50_reg_23218[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_66_fu_10171_p3 = ((or_ln346_13_reg_23223[0:0] == 1'b1) ? select_ln346_65_fu_10164_p3 : add_ln377_13_reg_23213);

assign select_ln346_67_fu_10205_p3 = ((and_ln895_51_fu_10199_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_68_fu_10219_p3 = ((xor_ln346_2_fu_10213_p2[0:0] == 1'b1) ? select_ln346_67_fu_10205_p3 : select_ln346_66_fu_10171_p3);

assign select_ln346_69_fu_10255_p3 = ((and_ln895_52_fu_10249_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_70_fu_10269_p3 = ((xor_ln346_3_fu_10263_p2[0:0] == 1'b1) ? select_ln346_69_fu_10255_p3 : select_ln346_68_fu_10219_p3);

assign select_ln346_71_fu_2722_p3 = ((and_ln895_53_fu_2686_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_72_fu_2730_p3 = ((or_ln346_14_fu_2716_p2[0:0] == 1'b1) ? select_ln346_71_fu_2722_p3 : add_ln377_14_fu_2586_p2);

assign select_ln346_73_fu_4058_p3 = ((and_ln895_54_reg_22584[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_74_fu_4065_p3 = ((or_ln346_15_fu_4053_p2[0:0] == 1'b1) ? select_ln346_73_fu_4058_p3 : add_ln377_15_reg_22569);

assign select_ln346_75_fu_4912_p3 = ((and_ln895_55_reg_22678[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_76_fu_4919_p3 = ((or_ln346_16_reg_22683[0:0] == 1'b1) ? select_ln346_75_fu_4912_p3 : add_ln377_16_reg_22673);

assign select_ln346_77_fu_5508_p3 = ((and_ln895_56_reg_22724[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_78_fu_5515_p3 = ((or_ln346_17_reg_22729[0:0] == 1'b1) ? select_ln346_77_fu_5508_p3 : add_ln377_17_reg_22719);

assign select_ln346_79_fu_5549_p3 = ((and_ln895_57_fu_5543_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_80_fu_5563_p3 = ((xor_ln346_4_fu_5557_p2[0:0] == 1'b1) ? select_ln346_79_fu_5549_p3 : select_ln346_78_fu_5515_p3);

assign select_ln346_81_fu_5605_p3 = ((and_ln895_58_fu_5593_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_82_fu_5613_p3 = ((xor_ln346_5_fu_5599_p2[0:0] == 1'b1) ? select_ln346_81_fu_5605_p3 : select_ln346_80_fu_5563_p3);

assign select_ln346_83_fu_6215_p3 = ((and_ln895_59_reg_22813[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_84_fu_6222_p3 = ((or_ln346_18_fu_6210_p2[0:0] == 1'b1) ? select_ln346_83_fu_6215_p3 : add_ln377_18_reg_22798);

assign select_ln346_85_fu_6887_p3 = ((and_ln895_60_reg_22912[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_86_fu_6894_p3 = ((or_ln346_19_reg_22917[0:0] == 1'b1) ? select_ln346_85_fu_6887_p3 : add_ln377_19_reg_22907);

assign select_ln346_87_fu_7093_p3 = ((and_ln895_61_fu_7057_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_88_fu_7101_p3 = ((or_ln346_20_fu_7087_p2[0:0] == 1'b1) ? select_ln346_87_fu_7093_p3 : add_ln377_20_fu_6955_p2);

assign select_ln346_89_fu_8369_p3 = ((and_ln895_62_reg_23013[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_90_fu_8376_p3 = ((or_ln346_21_reg_23018[0:0] == 1'b1) ? select_ln346_89_fu_8369_p3 : add_ln377_21_reg_23008);

assign select_ln346_91_fu_8416_p3 = ((and_ln895_63_fu_8404_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_92_fu_8424_p3 = ((xor_ln346_6_fu_8410_p2[0:0] == 1'b1) ? select_ln346_91_fu_8416_p3 : select_ln346_90_fu_8376_p3);

assign select_ln346_93_fu_8999_p3 = ((and_ln895_64_reg_23089[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_94_fu_9006_p3 = ((or_ln346_22_reg_23094[0:0] == 1'b1) ? select_ln346_93_fu_8999_p3 : add_ln377_22_reg_23084);

assign select_ln346_95_fu_9040_p3 = ((and_ln895_65_fu_9034_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_96_fu_9054_p3 = ((xor_ln346_7_fu_9048_p2[0:0] == 1'b1) ? select_ln346_95_fu_9040_p3 : select_ln346_94_fu_9006_p3);

assign select_ln346_97_fu_9096_p3 = ((and_ln895_66_fu_9084_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_98_fu_9104_p3 = ((xor_ln346_8_fu_9090_p2[0:0] == 1'b1) ? select_ln346_97_fu_9096_p3 : select_ln346_96_fu_9054_p3);

assign select_ln346_99_fu_9492_p3 = ((and_ln895_67_reg_23130[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln346_fu_1363_p3 = ((and_ln895_fu_1351_p2[0:0] == 1'b1) ? 21'd1048575 : 21'd1048576);

assign select_ln49_10_fu_19585_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_10_fu_19581_p1 : 20'd0);

assign select_ln49_11_fu_19602_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_11_fu_19598_p1 : 20'd0);

assign select_ln49_12_fu_19761_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_12_fu_19757_p1 : 20'd0);

assign select_ln49_13_fu_19778_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_13_fu_19774_p1 : 20'd0);

assign select_ln49_14_fu_19937_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_14_fu_19933_p1 : 20'd0);

assign select_ln49_15_fu_19954_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_15_fu_19950_p1 : 20'd0);

assign select_ln49_16_fu_20113_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_16_fu_20109_p1 : 20'd0);

assign select_ln49_17_fu_20130_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_17_fu_20126_p1 : 20'd0);

assign select_ln49_1_fu_18722_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_1_fu_18718_p1 : 20'd0);

assign select_ln49_2_fu_18881_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_2_fu_18877_p1 : 20'd0);

assign select_ln49_3_fu_18898_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_3_fu_18894_p1 : 20'd0);

assign select_ln49_4_fu_19057_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_4_fu_19053_p1 : 20'd0);

assign select_ln49_5_fu_19074_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_5_fu_19070_p1 : 20'd0);

assign select_ln49_6_fu_19233_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_6_fu_19229_p1 : 20'd0);

assign select_ln49_7_fu_19250_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_7_fu_19246_p1 : 20'd0);

assign select_ln49_8_fu_19409_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_8_fu_19405_p1 : 20'd0);

assign select_ln49_9_fu_19426_p3 = ((grp_fu_1194_p2[0:0] == 1'b1) ? trunc_ln1649_9_fu_19422_p1 : 20'd0);

assign select_ln49_fu_18705_p3 = ((grp_fu_1188_p2[0:0] == 1'b1) ? trunc_ln1649_fu_18701_p1 : 20'd0);

assign sext_ln1273_12_fu_2544_p1 = $signed(select_ln302_8_fu_2240_p3);

assign sext_ln1273_14_fu_8141_p1 = $signed(shl_ln1273_2_fu_8134_p3);

assign sext_ln1273_15_fu_8152_p1 = $signed(shl_ln1273_3_fu_8145_p3);

assign sext_ln1273_16_fu_3286_p1 = select_ln302_10_fu_2993_p3;

assign sext_ln1273_22_fu_4891_p1 = $signed(shl_ln1273_4_fu_4884_p3);

assign sext_ln1273_23_fu_4902_p1 = $signed(shl_ln1273_5_fu_4895_p3);

assign sext_ln1273_24_fu_7599_p1 = $signed(shl_ln1273_6_fu_7592_p3);

assign sext_ln1273_25_fu_7610_p1 = $signed(shl_ln1273_7_fu_7603_p3);

assign sext_ln1273_2_fu_1597_p1 = $signed(select_ln302_2_fu_1519_p3);

assign sext_ln1273_33_fu_10904_p1 = select_ln302_22_reg_23155;

assign sext_ln1273_37_fu_8721_p1 = select_ln302_23_fu_8709_p3;

assign sext_ln1273_38_fu_8733_p1 = $signed(shl_ln1273_8_fu_8725_p3);

assign sext_ln1273_39_fu_11359_p1 = $signed(shl_ln1273_9_fu_11352_p3);

assign sext_ln1273_40_fu_12212_p1 = select_ln346_139_fu_12187_p3;

assign sext_ln1273_41_fu_12216_p1 = select_ln346_139_fu_12187_p3;

assign sext_ln1273_42_fu_12220_p1 = select_ln346_139_fu_12187_p3;

assign sext_ln1273_43_fu_12224_p1 = select_ln346_139_fu_12187_p3;

assign sext_ln1273_44_fu_12228_p1 = select_ln346_139_fu_12187_p3;

assign sext_ln1273_45_fu_12232_p1 = select_ln346_145_fu_12206_p3;

assign sext_ln1273_46_fu_12537_p1 = select_ln346_145_reg_23375;

assign sext_ln1273_47_fu_12236_p1 = select_ln346_145_fu_12206_p3;

assign sext_ln1273_48_fu_12540_p1 = select_ln346_151_fu_12531_p3;

assign sext_ln1273_49_fu_12544_p1 = select_ln346_151_fu_12531_p3;

assign sext_ln1273_4_fu_3797_p1 = $signed(shl_ln1_fu_3790_p3);

assign sext_ln1273_50_fu_12638_p1 = $signed(shl_ln1273_11_fu_12631_p3);

assign sext_ln1273_5_fu_3808_p1 = $signed(shl_ln1273_1_fu_3801_p3);

assign sext_ln1273_6_fu_1601_p1 = select_ln302_19_fu_1589_p3;

assign sext_ln1347_10_fu_6679_p1 = mul_ln1273_6_reg_22657;

assign sext_ln1347_11_fu_6682_p1 = mul_ln1273_6_reg_22657;

assign sext_ln1347_12_fu_7395_p1 = mul_ln1273_7_reg_22703;

assign sext_ln1347_13_fu_8173_p1 = sub_ln1273_1_fu_8156_p2;

assign sext_ln1347_14_fu_8177_p1 = sub_ln1273_1_fu_8156_p2;

assign sext_ln1347_15_fu_8798_p1 = mul_ln1273_8_reg_22766;

assign sext_ln1347_16_fu_8801_p1 = mul_ln1273_8_reg_22766;

assign sext_ln1347_17_fu_9307_p1 = mul_ln1273_9_reg_22777;

assign sext_ln1347_18_fu_9310_p1 = mul_ln1273_9_reg_22777;

assign sext_ln1347_19_fu_3313_p1 = grp_fu_21456_p2;

assign sext_ln1347_1_fu_2332_p1 = mul_ln1273_1_reg_22425;

assign sext_ln1347_20_fu_3316_p1 = grp_fu_21456_p2;

assign sext_ln1347_21_fu_4084_p1 = mul_ln1273_14_reg_22500;

assign sext_ln1347_22_fu_4937_p1 = sub_ln1273_2_fu_4906_p2;

assign sext_ln1347_23_fu_4941_p1 = sub_ln1273_2_fu_4906_p2;

assign sext_ln1347_24_fu_5633_p1 = mul_ln1273_15_reg_22734;

assign sext_ln1347_25_fu_6241_p1 = mul_ln1273_16_reg_22745;

assign sext_ln1347_26_fu_6244_p1 = mul_ln1273_16_reg_22745;

assign sext_ln1347_27_fu_6912_p1 = mul_ln1273_17_reg_22824;

assign sext_ln1347_28_fu_7631_p1 = sub_ln1273_3_fu_7614_p2;

assign sext_ln1347_29_fu_7635_p1 = sub_ln1273_3_fu_7614_p2;

assign sext_ln1347_2_fu_3082_p1 = mul_ln1273_2_reg_22457;

assign sext_ln1347_30_fu_3487_p1 = grp_fu_21465_p2;

assign sext_ln1347_31_fu_3490_p1 = grp_fu_21465_p2;

assign sext_ln1347_32_fu_5806_p1 = grp_fu_21530_p2;

assign sext_ln1347_33_fu_6483_p1 = mul_ln1273_23_reg_22876;

assign sext_ln1347_34_fu_6486_p1 = mul_ln1273_23_reg_22876;

assign sext_ln1347_35_fu_10918_p1 = mul_ln1273_27_reg_23243;

assign sext_ln1347_36_fu_10921_p1 = mul_ln1273_27_reg_23243;

assign sext_ln1347_37_fu_11593_p1 = mul_ln1273_28_reg_23191;

assign sext_ln1347_38_fu_11596_p1 = mul_ln1273_28_reg_23191;

assign sext_ln1347_39_fu_11148_p1 = mul_ln1273_30_reg_23254;

assign sext_ln1347_3_fu_3829_p1 = sub_ln1273_fu_3812_p2;

assign sext_ln1347_40_fu_11151_p1 = mul_ln1273_30_reg_23254;

assign sext_ln1347_41_fu_11789_p1 = sub_ln1273_4_reg_23109;

assign sext_ln1347_42_fu_11792_p1 = sub_ln1273_4_reg_23109;

assign sext_ln1347_43_fu_11395_p1 = sub_ln1273_5_fu_11363_p2;

assign sext_ln1347_44_fu_11399_p1 = sub_ln1273_5_fu_11363_p2;

assign sext_ln1347_45_fu_11999_p1 = mul_ln1273_32_reg_23202;

assign sext_ln1347_46_fu_15174_p1 = grp_fu_21802_p2;

assign sext_ln1347_47_fu_15362_p1 = grp_fu_21810_p2;

assign sext_ln1347_48_fu_15365_p1 = grp_fu_21810_p2;

assign sext_ln1347_49_fu_15536_p1 = mul_ln1273_40_reg_23500;

assign sext_ln1347_4_fu_3833_p1 = sub_ln1273_fu_3812_p2;

assign sext_ln1347_50_fu_17322_p1 = mul_ln1273_41_reg_23676;

assign sext_ln1347_51_fu_15769_p1 = mul_ln1273_43_reg_23531;

assign sext_ln1347_52_fu_15772_p1 = mul_ln1273_43_reg_23531;

assign sext_ln1347_53_fu_17530_p1 = mul_ln1273_44_reg_23692;

assign sext_ln1347_54_fu_17533_p1 = mul_ln1273_44_reg_23692;

assign sext_ln1347_55_fu_16332_p1 = grp_fu_21855_p2;

assign sext_ln1347_56_fu_16520_p1 = grp_fu_21863_p2;

assign sext_ln1347_57_fu_16523_p1 = grp_fu_21863_p2;

assign sext_ln1347_58_fu_16694_p1 = mul_ln1273_52_reg_23562;

assign sext_ln1347_59_fu_18150_p1 = mul_ln1273_53_reg_23810;

assign sext_ln1347_5_fu_4672_p1 = mul_ln1273_3_reg_22473;

assign sext_ln1347_60_fu_16927_p1 = mul_ln1273_55_reg_23593;

assign sext_ln1347_61_fu_16930_p1 = mul_ln1273_55_reg_23593;

assign sext_ln1347_62_fu_18358_p1 = mul_ln1273_56_reg_23826;

assign sext_ln1347_63_fu_18361_p1 = mul_ln1273_56_reg_23826;

assign sext_ln1347_6_fu_4675_p1 = mul_ln1273_3_reg_22473;

assign sext_ln1347_7_fu_5293_p1 = mul_ln1273_4_reg_22527;

assign sext_ln1347_8_fu_5296_p1 = mul_ln1273_4_reg_22527;

assign sext_ln1347_9_fu_5987_p1 = mul_ln1273_5_reg_22646;

assign sext_ln1347_fu_2329_p1 = mul_ln1273_1_reg_22425;

assign sext_ln365_1_fu_10746_p1 = $signed(trunc_ln818_35_fu_10737_p4);

assign sext_ln365_2_fu_13297_p1 = $signed(trunc_ln818_39_fu_13288_p4);

assign sext_ln365_3_fu_13657_p1 = $signed(trunc_ln818_42_fu_13648_p4);

assign sext_ln365_4_fu_14028_p1 = $signed(trunc_ln818_47_fu_14019_p4);

assign sext_ln365_5_fu_16163_p1 = $signed(trunc_ln818_51_fu_16154_p4);

assign sext_ln365_6_fu_14395_p1 = $signed(trunc_ln818_54_fu_14386_p4);

assign sext_ln365_7_fu_14766_p1 = $signed(trunc_ln818_59_fu_14757_p4);

assign sext_ln365_fu_10572_p1 = $signed(trunc_ln818_32_fu_10563_p4);

assign sext_ln810_1_fu_12859_p1 = $signed(shl_ln1273_10_fu_12852_p3);

assign sext_ln810_fu_12848_p1 = $signed(shl_ln1273_s_fu_12841_p3);

assign sext_ln813_100_fu_10277_p1 = $signed(select_ln346_70_fu_10269_p3);

assign sext_ln813_101_fu_7980_p1 = $signed(shl_ln838_25_fu_7972_p3);

assign sext_ln813_102_fu_9555_p1 = $signed(select_ln346_102_fu_9547_p3);

assign sext_ln813_103_fu_8654_p1 = $signed(select_ln346_130_fu_8647_p3);

assign sext_ln813_104_fu_10914_p1 = shl_ln838_26_fu_10907_p3;

assign sext_ln813_105_fu_11589_p1 = shl_ln838_27_fu_11582_p3;

assign sext_ln813_106_fu_11144_p1 = shl_ln838_28_fu_11136_p3;

assign sext_ln813_107_fu_11785_p1 = shl_ln838_29_fu_11778_p3;

assign sext_ln813_108_fu_11391_p1 = shl_ln838_30_fu_11383_p3;

assign sext_ln813_109_fu_11995_p1 = shl_ln838_31_fu_11987_p3;

assign sext_ln813_110_fu_15170_p1 = shl_ln838_32_fu_15163_p3;

assign sext_ln813_111_fu_15358_p1 = shl_ln838_33_fu_15350_p3;

assign sext_ln813_112_fu_15532_p1 = shl_ln838_34_fu_15525_p3;

assign sext_ln813_113_fu_17318_p1 = shl_ln838_35_fu_17311_p3;

assign sext_ln813_114_fu_15765_p1 = shl_ln838_36_fu_15757_p3;

assign sext_ln813_115_fu_17526_p1 = shl_ln838_37_fu_17519_p3;

assign sext_ln813_116_fu_16328_p1 = shl_ln838_38_fu_16321_p3;

assign sext_ln813_117_fu_16516_p1 = shl_ln838_39_fu_16508_p3;

assign sext_ln813_118_fu_16690_p1 = shl_ln838_40_fu_16683_p3;

assign sext_ln813_119_fu_18146_p1 = shl_ln838_41_fu_18139_p3;

assign sext_ln813_120_fu_16923_p1 = shl_ln838_42_fu_16915_p3;

assign sext_ln813_121_fu_18354_p1 = shl_ln838_43_fu_18347_p3;

assign sext_ln813_122_fu_18559_p1 = reg_1200;

assign sext_ln813_123_fu_18563_p0 = Hxk_V_q1;

assign sext_ln813_123_fu_18563_p1 = sext_ln813_123_fu_18563_p0;

assign sext_ln813_124_fu_18630_p1 = reg_1204;

assign sext_ln813_125_fu_18634_p0 = Hxk_V_q0;

assign sext_ln813_125_fu_18634_p1 = sext_ln813_125_fu_18634_p0;

assign sext_ln813_126_fu_18735_p1 = reg_1208;

assign sext_ln813_127_fu_18739_p0 = Hxk_V_q1;

assign sext_ln813_127_fu_18739_p1 = sext_ln813_127_fu_18739_p0;

assign sext_ln813_128_fu_18806_p1 = reg_1212;

assign sext_ln813_129_fu_18810_p0 = Hxk_V_q0;

assign sext_ln813_129_fu_18810_p1 = sext_ln813_129_fu_18810_p0;

assign sext_ln813_130_fu_18911_p1 = reg_1216;

assign sext_ln813_131_fu_18915_p0 = Hxk_V_q1;

assign sext_ln813_131_fu_18915_p1 = sext_ln813_131_fu_18915_p0;

assign sext_ln813_132_fu_18982_p1 = reg_1220;

assign sext_ln813_133_fu_18986_p0 = Hxk_V_q0;

assign sext_ln813_133_fu_18986_p1 = sext_ln813_133_fu_18986_p0;

assign sext_ln813_134_fu_19087_p1 = reg_1224;

assign sext_ln813_135_fu_19091_p0 = Hxk_V_q1;

assign sext_ln813_135_fu_19091_p1 = sext_ln813_135_fu_19091_p0;

assign sext_ln813_136_fu_19158_p1 = reg_1228;

assign sext_ln813_137_fu_19162_p0 = Hxk_V_q0;

assign sext_ln813_137_fu_19162_p1 = sext_ln813_137_fu_19162_p0;

assign sext_ln813_138_fu_19263_p1 = reg_1232;

assign sext_ln813_139_fu_19267_p0 = Hxk_V_q1;

assign sext_ln813_139_fu_19267_p1 = sext_ln813_139_fu_19267_p0;

assign sext_ln813_140_fu_19334_p1 = reg_1236;

assign sext_ln813_141_fu_19338_p0 = Hxk_V_q0;

assign sext_ln813_141_fu_19338_p1 = sext_ln813_141_fu_19338_p0;

assign sext_ln813_142_fu_19439_p1 = reg_1240;

assign sext_ln813_143_fu_19443_p0 = Hxk_V_q1;

assign sext_ln813_143_fu_19443_p1 = sext_ln813_143_fu_19443_p0;

assign sext_ln813_144_fu_19510_p1 = reg_1244;

assign sext_ln813_145_fu_19514_p0 = Hxk_V_q0;

assign sext_ln813_145_fu_19514_p1 = sext_ln813_145_fu_19514_p0;

assign sext_ln813_146_fu_19615_p1 = reg_1248;

assign sext_ln813_147_fu_19619_p0 = Hxk_V_q1;

assign sext_ln813_147_fu_19619_p1 = sext_ln813_147_fu_19619_p0;

assign sext_ln813_148_fu_19686_p1 = reg_1252;

assign sext_ln813_149_fu_19690_p0 = Hxk_V_q0;

assign sext_ln813_149_fu_19690_p1 = sext_ln813_149_fu_19690_p0;

assign sext_ln813_150_fu_19791_p1 = reg_1256;

assign sext_ln813_151_fu_19795_p0 = Hxk_V_q1;

assign sext_ln813_151_fu_19795_p1 = sext_ln813_151_fu_19795_p0;

assign sext_ln813_152_fu_19862_p1 = reg_1260;

assign sext_ln813_153_fu_19866_p0 = Hxk_V_q0;

assign sext_ln813_153_fu_19866_p1 = sext_ln813_153_fu_19866_p0;

assign sext_ln813_154_fu_19967_p1 = reg_1264;

assign sext_ln813_155_fu_19971_p0 = Hxk_V_q1;

assign sext_ln813_155_fu_19971_p1 = sext_ln813_155_fu_19971_p0;

assign sext_ln813_156_fu_20038_p1 = reg_1268;

assign sext_ln813_157_fu_20042_p0 = Hxk_V_q0;

assign sext_ln813_157_fu_20042_p1 = sext_ln813_157_fu_20042_p0;

assign sext_ln813_158_fu_20143_p0 = temp7_q1;

assign sext_ln813_158_fu_20143_p1 = sext_ln813_158_fu_20143_p0;

assign sext_ln813_159_fu_20147_p1 = zk_admm_V_load_reg_23882;

assign sext_ln813_160_fu_20212_p0 = temp7_q0;

assign sext_ln813_160_fu_20212_p1 = sext_ln813_160_fu_20212_p0;

assign sext_ln813_161_fu_20216_p1 = zk_admm_V_load_1_reg_23888;

assign sext_ln813_162_fu_20281_p0 = temp7_q1;

assign sext_ln813_162_fu_20281_p1 = sext_ln813_162_fu_20281_p0;

assign sext_ln813_163_fu_20285_p1 = zk_admm_V_load_2_reg_23894;

assign sext_ln813_164_fu_20350_p0 = temp7_q0;

assign sext_ln813_164_fu_20350_p1 = sext_ln813_164_fu_20350_p0;

assign sext_ln813_165_fu_20354_p1 = zk_admm_V_load_3_reg_23900;

assign sext_ln813_166_fu_20419_p0 = temp7_q1;

assign sext_ln813_166_fu_20419_p1 = sext_ln813_166_fu_20419_p0;

assign sext_ln813_167_fu_20423_p1 = zk_admm_V_load_4_reg_23906;

assign sext_ln813_168_fu_20488_p0 = temp7_q0;

assign sext_ln813_168_fu_20488_p1 = sext_ln813_168_fu_20488_p0;

assign sext_ln813_169_fu_20492_p1 = zk_admm_V_load_5_reg_23912;

assign sext_ln813_170_fu_20557_p0 = temp7_q1;

assign sext_ln813_170_fu_20557_p1 = sext_ln813_170_fu_20557_p0;

assign sext_ln813_171_fu_20561_p1 = zk_admm_V_load_6_reg_23918;

assign sext_ln813_172_fu_20626_p0 = temp7_q0;

assign sext_ln813_172_fu_20626_p1 = sext_ln813_172_fu_20626_p0;

assign sext_ln813_173_fu_20630_p1 = zk_admm_V_load_7_reg_23924;

assign sext_ln813_174_fu_20695_p0 = temp7_q1;

assign sext_ln813_174_fu_20695_p1 = sext_ln813_174_fu_20695_p0;

assign sext_ln813_175_fu_20699_p1 = zk_admm_V_load_8_reg_23930;

assign sext_ln813_176_fu_20764_p0 = temp7_q0;

assign sext_ln813_176_fu_20764_p1 = sext_ln813_176_fu_20764_p0;

assign sext_ln813_177_fu_20768_p1 = zk_admm_V_load_9_reg_23936;

assign sext_ln813_178_fu_20833_p0 = temp7_q1;

assign sext_ln813_178_fu_20833_p1 = sext_ln813_178_fu_20833_p0;

assign sext_ln813_179_fu_20837_p1 = zk_admm_V_load_10_reg_23942;

assign sext_ln813_180_fu_20902_p0 = temp7_q0;

assign sext_ln813_180_fu_20902_p1 = sext_ln813_180_fu_20902_p0;

assign sext_ln813_181_fu_20906_p1 = zk_admm_V_load_11_reg_23948;

assign sext_ln813_182_fu_20971_p0 = temp7_q1;

assign sext_ln813_182_fu_20971_p1 = sext_ln813_182_fu_20971_p0;

assign sext_ln813_183_fu_20975_p1 = zk_admm_V_load_12_reg_23954;

assign sext_ln813_184_fu_21040_p0 = temp7_q0;

assign sext_ln813_184_fu_21040_p1 = sext_ln813_184_fu_21040_p0;

assign sext_ln813_185_fu_21044_p1 = zk_admm_V_load_13_reg_23960;

assign sext_ln813_186_fu_21109_p0 = temp7_q1;

assign sext_ln813_186_fu_21109_p1 = sext_ln813_186_fu_21109_p0;

assign sext_ln813_187_fu_21113_p1 = zk_admm_V_load_14_reg_23966;

assign sext_ln813_188_fu_21178_p0 = temp7_q0;

assign sext_ln813_188_fu_21178_p1 = sext_ln813_188_fu_21178_p0;

assign sext_ln813_189_fu_21182_p1 = zk_admm_V_load_15_reg_23972;

assign sext_ln813_190_fu_21247_p0 = temp7_q1;

assign sext_ln813_190_fu_21247_p1 = sext_ln813_190_fu_21247_p0;

assign sext_ln813_191_fu_21251_p1 = zk_admm_V_load_16_reg_23978;

assign sext_ln813_192_fu_21316_p0 = temp7_q0;

assign sext_ln813_192_fu_21316_p1 = sext_ln813_192_fu_21316_p0;

assign sext_ln813_193_fu_21320_p1 = zk_admm_V_load_17_reg_23984;

assign sext_ln813_36_fu_1313_p1 = reg_1200;

assign sext_ln813_37_fu_1379_p0 = temp_q0;

assign sext_ln813_37_fu_1379_p1 = sext_ln813_37_fu_1379_p0;

assign sext_ln813_38_fu_1383_p1 = reg_1204;

assign sext_ln813_39_fu_1457_p0 = temp_q1;

assign sext_ln813_39_fu_1457_p1 = sext_ln813_39_fu_1457_p0;

assign sext_ln813_40_fu_1461_p1 = reg_1208;

assign sext_ln813_41_fu_1609_p0 = temp_q1;

assign sext_ln813_41_fu_1609_p1 = sext_ln813_41_fu_1609_p0;

assign sext_ln813_42_fu_1613_p1 = reg_1216;

assign sext_ln813_43_fu_1527_p0 = temp_q0;

assign sext_ln813_43_fu_1527_p1 = sext_ln813_43_fu_1527_p0;

assign sext_ln813_44_fu_1531_p1 = reg_1212;

assign sext_ln813_45_fu_1679_p0 = temp_q0;

assign sext_ln813_45_fu_1679_p1 = sext_ln813_45_fu_1679_p0;

assign sext_ln813_46_fu_1683_p1 = reg_1220;

assign sext_ln813_47_fu_1837_p0 = temp_q1;

assign sext_ln813_47_fu_1837_p1 = sext_ln813_47_fu_1837_p0;

assign sext_ln813_48_fu_1841_p1 = reg_1224;

assign sext_ln813_49_fu_1907_p0 = temp_q0;

assign sext_ln813_49_fu_1907_p1 = sext_ln813_49_fu_1907_p0;

assign sext_ln813_50_fu_1911_p1 = reg_1228;

assign sext_ln813_51_fu_2178_p0 = temp_q1;

assign sext_ln813_51_fu_2178_p1 = sext_ln813_51_fu_2178_p0;

assign sext_ln813_52_fu_2182_p1 = reg_1232;

assign sext_ln813_53_fu_2248_p0 = temp_q0;

assign sext_ln813_53_fu_2248_p1 = sext_ln813_53_fu_2248_p0;

assign sext_ln813_54_fu_2252_p1 = reg_1236;

assign sext_ln813_55_fu_2931_p0 = temp_q1;

assign sext_ln813_55_fu_2931_p1 = sext_ln813_55_fu_2931_p0;

assign sext_ln813_56_fu_2935_p1 = reg_1240;

assign sext_ln813_57_fu_3001_p0 = temp_q0;

assign sext_ln813_57_fu_3001_p1 = sext_ln813_57_fu_3001_p0;

assign sext_ln813_58_fu_3005_p1 = reg_1244;

assign sext_ln813_59_fu_3650_p0 = temp_q1;

assign sext_ln813_59_fu_3650_p1 = sext_ln813_59_fu_3650_p0;

assign sext_ln813_60_fu_3654_p1 = reg_1248;

assign sext_ln813_61_fu_3720_p0 = temp_q0;

assign sext_ln813_61_fu_3720_p1 = sext_ln813_61_fu_3720_p0;

assign sext_ln813_62_fu_3724_p1 = reg_1252;

assign sext_ln813_63_fu_4507_p0 = temp_q1;

assign sext_ln813_63_fu_4507_p1 = sext_ln813_63_fu_4507_p0;

assign sext_ln813_64_fu_4511_p1 = reg_1256;

assign sext_ln813_65_fu_4577_p0 = temp_q0;

assign sext_ln813_65_fu_4577_p1 = sext_ln813_65_fu_4577_p0;

assign sext_ln813_66_fu_4581_p1 = reg_1260;

assign sext_ln813_67_fu_5142_p0 = temp_q1;

assign sext_ln813_67_fu_5142_p1 = sext_ln813_67_fu_5142_p0;

assign sext_ln813_68_fu_5146_p1 = reg_1264;

assign sext_ln813_69_fu_5212_p0 = temp_q0;

assign sext_ln813_69_fu_5212_p1 = sext_ln813_69_fu_5212_p0;

assign sext_ln813_70_fu_5216_p1 = reg_1268;

assign sext_ln813_71_fu_1272_p1 = $signed(p_read);

assign sext_ln813_72_fu_1276_p1 = $signed(p_read1);

assign sext_ln813_73_fu_1280_p1 = $signed(p_read2);

assign sext_ln813_74_fu_2325_p1 = shl_ln_fu_2318_p3;

assign sext_ln813_75_fu_3078_p1 = shl_ln838_1_fu_3071_p3;

assign sext_ln813_76_fu_3825_p1 = shl_ln838_2_fu_3818_p3;

assign sext_ln813_77_fu_4668_p1 = shl_ln838_3_fu_4660_p3;

assign sext_ln813_78_fu_5289_p1 = shl_ln838_4_fu_5282_p3;

assign sext_ln813_79_fu_5983_p1 = shl_ln838_5_fu_5976_p3;

assign sext_ln813_80_fu_6675_p1 = shl_ln838_6_fu_6668_p3;

assign sext_ln813_81_fu_7391_p1 = shl_ln838_7_fu_7384_p3;

assign sext_ln813_82_fu_8169_p1 = shl_ln838_8_fu_8162_p3;

assign sext_ln813_83_fu_8794_p1 = shl_ln838_9_fu_8786_p3;

assign sext_ln813_84_fu_9303_p1 = shl_ln838_s_fu_9296_p3;

assign sext_ln813_85_fu_9677_p1 = $signed(shl_ln838_10_fu_9669_p3);

assign sext_ln813_86_fu_9988_p1 = $signed(shl_ln838_11_fu_9980_p3);

assign sext_ln813_87_fu_3309_p1 = shl_ln838_12_fu_3302_p3;

assign sext_ln813_88_fu_4080_p1 = shl_ln838_13_fu_4072_p3;

assign sext_ln813_89_fu_4933_p1 = shl_ln838_14_fu_4925_p3;

assign sext_ln813_90_fu_5629_p1 = shl_ln838_15_fu_5621_p3;

assign sext_ln813_91_fu_6237_p1 = shl_ln838_16_fu_6229_p3;

assign sext_ln813_92_fu_6908_p1 = shl_ln838_17_fu_6900_p3;

assign sext_ln813_93_fu_7627_p1 = shl_ln838_18_fu_7620_p3;

assign sext_ln813_94_fu_8440_p1 = $signed(shl_ln838_19_fu_8432_p3);

assign sext_ln813_95_fu_9120_p1 = $signed(shl_ln838_20_fu_9112_p3);

assign sext_ln813_96_fu_3483_p1 = shl_ln838_21_fu_3476_p3;

assign sext_ln813_97_fu_5802_p1 = shl_ln838_22_fu_5795_p3;

assign sext_ln813_98_fu_6479_p1 = shl_ln838_23_fu_6471_p3;

assign sext_ln813_99_fu_7230_p1 = $signed(shl_ln838_24_fu_7222_p3);

assign sext_ln813_fu_1309_p0 = temp_q1;

assign sext_ln813_fu_1309_p1 = sext_ln813_fu_1309_p0;

assign sext_ln818_1_fu_13831_p1 = $signed(trunc_ln818_44_fu_13822_p4);

assign sext_ln818_2_fu_14569_p1 = $signed(trunc_ln818_56_fu_14560_p4);

assign sext_ln818_fu_10382_p1 = $signed(trunc_ln818_29_fu_10373_p4);

assign sext_ln856_1_fu_11349_p1 = add_ln377_36_reg_23285;

assign sext_ln856_2_fu_15045_p1 = add_ln377_40_reg_23465;

assign sext_ln856_3_fu_15333_p1 = add_ln377_43_reg_23485;

assign sext_ln856_4_fu_15740_p1 = add_ln377_48_reg_23516;

assign sext_ln856_5_fu_17845_p1 = add_ln377_52_reg_23723;

assign sext_ln856_6_fu_16491_p1 = add_ln377_55_reg_23547;

assign sext_ln856_7_fu_16898_p1 = add_ln377_60_reg_23578;

assign sext_ln856_fu_11119_p1 = add_ln377_33_reg_23270;

assign shl_ln1273_10_fu_12852_p3 = {{select_ln346_151_reg_23427}, {14'd0}};

assign shl_ln1273_11_fu_12631_p3 = {{select_ln346_139_reg_23370}, {14'd0}};

assign shl_ln1273_1_fu_3801_p3 = {{select_ln302_3_reg_22388}, {5'd0}};

assign shl_ln1273_2_fu_8134_p3 = {{select_ln302_9_reg_22451}, {7'd0}};

assign shl_ln1273_3_fu_8145_p3 = {{select_ln302_9_reg_22451}, {5'd0}};

assign shl_ln1273_4_fu_4884_p3 = {{select_ln302_5_reg_22394}, {7'd0}};

assign shl_ln1273_5_fu_4895_p3 = {{select_ln302_5_reg_22394}, {5'd0}};

assign shl_ln1273_6_fu_7592_p3 = {{select_ln302_11_reg_22516}, {7'd0}};

assign shl_ln1273_7_fu_7603_p3 = {{select_ln302_11_reg_22516}, {5'd0}};

assign shl_ln1273_8_fu_8725_p3 = {{select_ln302_23_fu_8709_p3}, {8'd0}};

assign shl_ln1273_9_fu_11352_p3 = {{select_ln302_22_reg_23155}, {8'd0}};

assign shl_ln1273_s_fu_12841_p3 = {{select_ln346_145_reg_23375}, {14'd0}};

assign shl_ln1_fu_3790_p3 = {{select_ln302_3_reg_22388}, {7'd0}};

assign shl_ln838_10_fu_9669_p3 = {{select_ln346_58_fu_9663_p3}, {14'd0}};

assign shl_ln838_11_fu_9980_p3 = {{select_ln346_64_fu_9972_p3}, {14'd0}};

assign shl_ln838_12_fu_3302_p3 = {{select_ln346_72_reg_22495}, {14'd0}};

assign shl_ln838_13_fu_4072_p3 = {{select_ln346_74_fu_4065_p3}, {14'd0}};

assign shl_ln838_14_fu_4925_p3 = {{select_ln346_76_fu_4919_p3}, {14'd0}};

assign shl_ln838_15_fu_5621_p3 = {{select_ln346_82_fu_5613_p3}, {14'd0}};

assign shl_ln838_16_fu_6229_p3 = {{select_ln346_84_fu_6222_p3}, {14'd0}};

assign shl_ln838_17_fu_6900_p3 = {{select_ln346_86_fu_6894_p3}, {14'd0}};

assign shl_ln838_18_fu_7620_p3 = {{select_ln346_88_reg_22962}, {14'd0}};

assign shl_ln838_19_fu_8432_p3 = {{select_ln346_92_fu_8424_p3}, {14'd0}};

assign shl_ln838_1_fu_3071_p3 = {{select_ln346_38_reg_22463}, {14'd0}};

assign shl_ln838_20_fu_9112_p3 = {{select_ln346_98_fu_9104_p3}, {14'd0}};

assign shl_ln838_21_fu_3476_p3 = {{select_ln346_104_reg_22511}, {14'd0}};

assign shl_ln838_22_fu_5795_p3 = {{select_ln346_114_reg_22693}, {14'd0}};

assign shl_ln838_23_fu_6471_p3 = {{select_ln346_116_fu_6464_p3}, {14'd0}};

assign shl_ln838_24_fu_7222_p3 = {{select_ln346_122_fu_7214_p3}, {14'd0}};

assign shl_ln838_25_fu_7972_p3 = {{select_ln346_128_fu_7964_p3}, {14'd0}};

assign shl_ln838_26_fu_10907_p3 = {{select_ln346_135_reg_23265}, {14'd0}};

assign shl_ln838_27_fu_11582_p3 = {{select_ln346_137_reg_23300}, {14'd0}};

assign shl_ln838_28_fu_11136_p3 = {{select_ln346_141_fu_11129_p3}, {14'd0}};

assign shl_ln838_29_fu_11778_p3 = {{select_ln346_143_reg_23305}, {14'd0}};

assign shl_ln838_2_fu_3818_p3 = {{select_ln346_40_reg_22522}, {14'd0}};

assign shl_ln838_30_fu_11383_p3 = {{select_ln346_147_fu_11376_p3}, {14'd0}};

assign shl_ln838_31_fu_11987_p3 = {{select_ln346_149_fu_11981_p3}, {14'd0}};

assign shl_ln838_32_fu_15163_p3 = {{select_ln346_165_reg_23480}, {14'd0}};

assign shl_ln838_33_fu_15350_p3 = {{select_ln346_171_fu_15343_p3}, {14'd0}};

assign shl_ln838_34_fu_15525_p3 = {{select_ln346_177_reg_23506}, {14'd0}};

assign shl_ln838_35_fu_17311_p3 = {{select_ln346_179_reg_23682}, {14'd0}};

assign shl_ln838_36_fu_15757_p3 = {{select_ln346_183_fu_15750_p3}, {14'd0}};

assign shl_ln838_37_fu_17519_p3 = {{select_ln346_185_reg_23698}, {14'd0}};

assign shl_ln838_38_fu_16321_p3 = {{select_ln346_201_reg_23542}, {14'd0}};

assign shl_ln838_39_fu_16508_p3 = {{select_ln346_207_fu_16501_p3}, {14'd0}};

assign shl_ln838_3_fu_4660_p3 = {{select_ln346_42_fu_4654_p3}, {14'd0}};

assign shl_ln838_40_fu_16683_p3 = {{select_ln346_213_reg_23568}, {14'd0}};

assign shl_ln838_41_fu_18139_p3 = {{select_ln346_215_reg_23816}, {14'd0}};

assign shl_ln838_42_fu_16915_p3 = {{select_ln346_219_fu_16908_p3}, {14'd0}};

assign shl_ln838_43_fu_18347_p3 = {{select_ln346_221_reg_23832}, {14'd0}};

assign shl_ln838_4_fu_5282_p3 = {{select_ln346_44_reg_22698}, {14'd0}};

assign shl_ln838_5_fu_5976_p3 = {{select_ln346_46_reg_22761}, {14'd0}};

assign shl_ln838_6_fu_6668_p3 = {{select_ln346_48_reg_22892}, {14'd0}};

assign shl_ln838_7_fu_7384_p3 = {{select_ln346_50_reg_22947}, {14'd0}};

assign shl_ln838_8_fu_8162_p3 = {{select_ln346_52_reg_23003}, {14'd0}};

assign shl_ln838_9_fu_8786_p3 = {{select_ln346_54_fu_8780_p3}, {14'd0}};

assign shl_ln838_s_fu_9296_p3 = {{select_ln346_56_reg_23120}, {14'd0}};

assign shl_ln_fu_2318_p3 = {{select_ln346_36_reg_22431}, {14'd0}};

assign sub_ln1273_1_fu_8156_p2 = ($signed(sext_ln1273_14_fu_8141_p1) - $signed(sext_ln1273_15_fu_8152_p1));

assign sub_ln1273_2_fu_4906_p2 = ($signed(sext_ln1273_23_fu_4902_p1) - $signed(sext_ln1273_22_fu_4891_p1));

assign sub_ln1273_3_fu_7614_p2 = ($signed(sext_ln1273_24_fu_7599_p1) - $signed(sext_ln1273_25_fu_7610_p1));

assign sub_ln1273_4_fu_8753_p2 = ($signed(sext_ln1273_37_fu_8721_p1) - $signed(sext_ln1273_38_fu_8733_p1));

assign sub_ln1273_5_fu_11363_p2 = ($signed(sext_ln1273_33_fu_10904_p1) - $signed(sext_ln1273_39_fu_11359_p1));

assign sub_ln1273_6_fu_12642_p2 = ($signed(36'd0) - $signed(sext_ln1273_50_fu_12638_p1));

assign sub_ln1273_7_fu_12863_p2 = ($signed(36'd0) - $signed(sext_ln810_fu_12848_p1));

assign sub_ln1273_8_fu_13012_p2 = ($signed(36'd0) - $signed(sext_ln810_1_fu_12859_p1));

assign sub_ln1273_fu_3812_p2 = ($signed(sext_ln1273_5_fu_3808_p1) - $signed(sext_ln1273_4_fu_3797_p1));

assign sub_ln1347_1_fu_1823_p2 = (trunc_ln1273_3_fu_1815_p3 - trunc_ln1273_2_fu_1803_p3);

assign sub_ln1347_2_fu_8759_p2 = (trunc_ln1273_10_fu_8749_p1 - trunc_ln1273_4_fu_8741_p3);

assign sub_ln1347_3_fu_9642_p2 = (trunc_ln1273_12_fu_9638_p1 - trunc_ln1273_5_fu_9630_p3);

assign sub_ln1347_fu_1777_p2 = (trunc_ln1273_1_fu_1769_p3 - trunc_ln2_fu_1757_p3);

assign sub_ln1348_18_fu_9559_p2 = ($signed(sext_ln813_102_fu_9555_p1) - $signed(sext_ln813_72_reg_21988));

assign sub_ln1348_19_fu_8658_p2 = ($signed(sext_ln813_103_fu_8654_p1) - $signed(sext_ln813_73_reg_21993));

assign sub_ln1348_fu_10281_p2 = ($signed(sext_ln813_100_fu_10277_p1) - $signed(sext_ln813_71_reg_21983));

assign tmp_100_fu_4771_p3 = add_ln1347_21_fu_4678_p2[32'd35];

assign tmp_101_fu_5311_p3 = add_ln1347_22_fu_5299_p2[32'd35];

assign tmp_102_fu_5329_p3 = add_ln810_4_fu_5305_p2[32'd34];

assign tmp_104_fu_5346_p3 = add_ln377_5_fu_5340_p2[32'd20];

assign tmp_105_fu_5366_p3 = add_ln1347_22_fu_5299_p2[32'd35];

assign tmp_106_fu_5392_p3 = add_ln1347_22_fu_5299_p2[32'd35];

assign tmp_107_fu_6001_p3 = add_ln1347_23_fu_5990_p2[32'd35];

assign tmp_108_fu_6019_p3 = add_ln810_5_fu_5996_p2[32'd34];

assign tmp_110_fu_6036_p3 = add_ln377_6_fu_6030_p2[32'd20];

assign tmp_111_fu_6056_p3 = add_ln1347_23_fu_5990_p2[32'd35];

assign tmp_112_fu_6082_p3 = add_ln1347_23_fu_5990_p2[32'd35];

assign tmp_113_fu_6697_p3 = add_ln1347_24_fu_6685_p2[32'd35];

assign tmp_114_fu_6715_p3 = add_ln810_6_fu_6691_p2[32'd34];

assign tmp_116_fu_6732_p3 = add_ln377_7_fu_6726_p2[32'd20];

assign tmp_117_fu_6752_p3 = add_ln1347_24_fu_6685_p2[32'd35];

assign tmp_118_fu_6778_p3 = add_ln1347_24_fu_6685_p2[32'd35];

assign tmp_119_fu_7409_p3 = add_ln1347_25_fu_7398_p2[32'd35];

assign tmp_120_fu_7427_p3 = add_ln810_7_fu_7404_p2[32'd34];

assign tmp_122_fu_7444_p3 = add_ln377_8_fu_7438_p2[32'd20];

assign tmp_123_fu_7464_p3 = add_ln1347_25_fu_7398_p2[32'd35];

assign tmp_124_fu_7490_p3 = add_ln1347_25_fu_7398_p2[32'd35];

assign tmp_125_fu_8193_p3 = add_ln1347_26_fu_8181_p2[32'd35];

assign tmp_126_fu_8211_p3 = add_ln810_8_fu_8187_p2[32'd34];

assign tmp_127_fu_8219_p3 = sub_ln1273_1_fu_8156_p2[32'd13];

assign tmp_128_fu_8237_p3 = add_ln377_9_fu_8231_p2[32'd20];

assign tmp_129_fu_8257_p3 = add_ln1347_26_fu_8181_p2[32'd35];

assign tmp_130_fu_8283_p3 = add_ln1347_26_fu_8181_p2[32'd35];

assign tmp_131_fu_8816_p3 = add_ln1347_27_fu_8804_p2[32'd35];

assign tmp_132_fu_8834_p3 = add_ln810_9_fu_8810_p2[32'd34];

assign tmp_134_fu_8851_p3 = add_ln377_10_fu_8845_p2[32'd20];

assign tmp_135_fu_8871_p3 = add_ln1347_27_fu_8804_p2[32'd35];

assign tmp_136_fu_8897_p3 = add_ln1347_27_fu_8804_p2[32'd35];

assign tmp_137_fu_9325_p3 = add_ln1347_28_fu_9313_p2[32'd35];

assign tmp_138_fu_9343_p3 = add_ln810_10_fu_9319_p2[32'd34];

assign tmp_140_fu_9360_p3 = add_ln377_11_fu_9354_p2[32'd20];

assign tmp_141_fu_9380_p3 = add_ln1347_28_fu_9313_p2[32'd35];

assign tmp_142_fu_9406_p3 = add_ln1347_28_fu_9313_p2[32'd35];

assign tmp_143_fu_9686_p3 = add_ln1347_29_fu_9681_p2[32'd35];

assign tmp_144_fu_9704_p3 = add_ln1347_29_fu_9681_p2[32'd34];

assign tmp_146_fu_9721_p3 = add_ln377_12_fu_9715_p2[32'd20];

assign tmp_147_fu_9741_p3 = add_ln1347_29_fu_9681_p2[32'd35];

assign tmp_148_fu_9767_p3 = add_ln1347_29_fu_9681_p2[32'd35];

assign tmp_149_fu_9880_p3 = select_ln346_60_fu_9874_p3[32'd20];

assign tmp_150_fu_9888_p3 = select_ln346_60_fu_9874_p3[32'd20];

assign tmp_151_fu_9930_p3 = select_ln346_62_fu_9922_p3[32'd20];

assign tmp_152_fu_9938_p3 = select_ln346_62_fu_9922_p3[32'd20];

assign tmp_153_fu_9997_p3 = add_ln1347_30_fu_9992_p2[32'd35];

assign tmp_154_fu_10015_p3 = add_ln1347_30_fu_9992_p2[32'd34];

assign tmp_156_fu_10032_p3 = add_ln377_13_fu_10026_p2[32'd20];

assign tmp_157_fu_10052_p3 = add_ln1347_30_fu_9992_p2[32'd35];

assign tmp_158_fu_10078_p3 = add_ln1347_30_fu_9992_p2[32'd35];

assign tmp_159_fu_10177_p3 = select_ln346_66_fu_10171_p3[32'd20];

assign tmp_160_fu_10185_p3 = select_ln346_66_fu_10171_p3[32'd20];

assign tmp_161_fu_10227_p3 = select_ln346_68_fu_10219_p3[32'd20];

assign tmp_162_fu_10235_p3 = select_ln346_68_fu_10219_p3[32'd20];

assign tmp_163_fu_2552_p3 = grp_fu_21418_p2[32'd34];

assign tmp_164_fu_2568_p3 = grp_fu_21418_p2[32'd34];

assign tmp_165_fu_2575_p3 = grp_fu_21418_p2[32'd13];

assign tmp_166_fu_2592_p3 = add_ln377_14_fu_2586_p2[32'd20];

assign tmp_167_fu_2612_p3 = grp_fu_21418_p2[32'd34];

assign tmp_168_fu_2637_p3 = grp_fu_21418_p2[32'd34];

assign tmp_169_fu_3331_p3 = add_ln1347_31_fu_3319_p2[32'd35];

assign tmp_170_fu_3349_p3 = add_ln810_11_fu_3325_p2[32'd34];

assign tmp_171_fu_3357_p3 = grp_fu_21456_p2[32'd13];

assign tmp_172_fu_3374_p3 = add_ln377_15_fu_3368_p2[32'd20];

assign tmp_173_fu_3388_p3 = add_ln1347_31_fu_3319_p2[32'd35];

assign tmp_174_fu_3414_p3 = add_ln1347_31_fu_3319_p2[32'd35];

assign tmp_175_fu_4098_p3 = add_ln1347_32_fu_4087_p2[32'd35];

assign tmp_176_fu_4116_p3 = add_ln810_12_fu_4093_p2[32'd34];

assign tmp_178_fu_4133_p3 = add_ln377_16_fu_4127_p2[32'd20];

assign tmp_179_fu_4153_p3 = add_ln1347_32_fu_4087_p2[32'd35];

assign tmp_180_fu_4179_p3 = add_ln1347_32_fu_4087_p2[32'd35];

assign tmp_181_fu_4957_p3 = add_ln1347_33_fu_4945_p2[32'd35];

assign tmp_182_fu_4975_p3 = add_ln810_13_fu_4951_p2[32'd34];

assign tmp_184_fu_4992_p3 = add_ln377_17_fu_4986_p2[32'd20];

assign tmp_185_fu_5012_p3 = add_ln1347_33_fu_4945_p2[32'd35];

assign tmp_186_fu_5038_p3 = add_ln1347_33_fu_4945_p2[32'd35];

assign tmp_187_fu_5521_p3 = select_ln346_78_fu_5515_p3[32'd20];

assign tmp_188_fu_5529_p3 = select_ln346_78_fu_5515_p3[32'd20];

assign tmp_189_fu_5571_p3 = select_ln346_80_fu_5563_p3[32'd20];

assign tmp_190_fu_5579_p3 = select_ln346_80_fu_5563_p3[32'd20];

assign tmp_191_fu_5647_p3 = add_ln1347_34_fu_5636_p2[32'd35];

assign tmp_192_fu_5665_p3 = add_ln810_14_fu_5642_p2[32'd34];

assign tmp_194_fu_5682_p3 = add_ln377_18_fu_5676_p2[32'd20];

assign tmp_195_fu_5696_p3 = add_ln1347_34_fu_5636_p2[32'd35];

assign tmp_196_fu_5722_p3 = add_ln1347_34_fu_5636_p2[32'd35];

assign tmp_197_fu_6259_p3 = add_ln1347_35_fu_6247_p2[32'd35];

assign tmp_198_fu_6277_p3 = add_ln810_15_fu_6253_p2[32'd34];

assign tmp_200_fu_6294_p3 = add_ln377_19_fu_6288_p2[32'd20];

assign tmp_201_fu_6314_p3 = add_ln1347_35_fu_6247_p2[32'd35];

assign tmp_202_fu_6340_p3 = add_ln1347_35_fu_6247_p2[32'd35];

assign tmp_203_fu_6926_p3 = add_ln1347_36_fu_6915_p2[32'd35];

assign tmp_204_fu_6944_p3 = add_ln810_16_fu_6921_p2[32'd34];

assign tmp_206_fu_6961_p3 = add_ln377_20_fu_6955_p2[32'd20];

assign tmp_207_fu_6981_p3 = add_ln1347_36_fu_6915_p2[32'd35];

assign tmp_208_fu_7007_p3 = add_ln1347_36_fu_6915_p2[32'd35];

assign tmp_209_fu_7651_p3 = add_ln1347_37_fu_7639_p2[32'd35];

assign tmp_210_fu_7669_p3 = add_ln810_17_fu_7645_p2[32'd34];

assign tmp_211_fu_7677_p3 = sub_ln1273_3_fu_7614_p2[32'd13];

assign tmp_212_fu_7695_p3 = add_ln377_21_fu_7689_p2[32'd20];

assign tmp_213_fu_7715_p3 = add_ln1347_37_fu_7639_p2[32'd35];

assign tmp_214_fu_7741_p3 = add_ln1347_37_fu_7639_p2[32'd35];

assign tmp_215_fu_8382_p3 = select_ln346_90_fu_8376_p3[32'd20];

assign tmp_216_fu_8390_p3 = select_ln346_90_fu_8376_p3[32'd20];

assign tmp_217_fu_8449_p3 = add_ln1347_38_fu_8444_p2[32'd35];

assign tmp_218_fu_8467_p3 = add_ln1347_38_fu_8444_p2[32'd34];

assign tmp_220_fu_8484_p3 = add_ln377_22_fu_8478_p2[32'd20];

assign tmp_221_fu_8504_p3 = add_ln1347_38_fu_8444_p2[32'd35];

assign tmp_222_fu_8530_p3 = add_ln1347_38_fu_8444_p2[32'd35];

assign tmp_223_fu_9012_p3 = select_ln346_94_fu_9006_p3[32'd20];

assign tmp_224_fu_9020_p3 = select_ln346_94_fu_9006_p3[32'd20];

assign tmp_225_fu_9062_p3 = select_ln346_96_fu_9054_p3[32'd20];

assign tmp_226_fu_9070_p3 = select_ln346_96_fu_9054_p3[32'd20];

assign tmp_227_fu_9129_p3 = add_ln1347_39_fu_9124_p2[32'd35];

assign tmp_228_fu_9147_p3 = add_ln1347_39_fu_9124_p2[32'd34];

assign tmp_230_fu_9164_p3 = add_ln377_23_fu_9158_p2[32'd20];

assign tmp_231_fu_9184_p3 = add_ln1347_39_fu_9124_p2[32'd35];

assign tmp_232_fu_9210_p3 = add_ln1347_39_fu_9124_p2[32'd35];

assign tmp_233_fu_9505_p3 = select_ln346_100_fu_9499_p3[32'd20];

assign tmp_234_fu_9513_p3 = select_ln346_100_fu_9499_p3[32'd20];

assign tmp_235_fu_2745_p3 = grp_fu_21437_p2[32'd34];

assign tmp_236_fu_2761_p3 = grp_fu_21437_p2[32'd34];

assign tmp_237_fu_2768_p3 = grp_fu_21437_p2[32'd13];

assign tmp_238_fu_2785_p3 = add_ln377_24_fu_2779_p2[32'd20];

assign tmp_239_fu_2805_p3 = grp_fu_21437_p2[32'd34];

assign tmp_240_fu_2830_p3 = grp_fu_21437_p2[32'd34];

assign tmp_241_fu_3505_p3 = add_ln1347_40_fu_3493_p2[32'd35];

assign tmp_242_fu_3523_p3 = add_ln810_18_fu_3499_p2[32'd34];

assign tmp_243_fu_3531_p3 = grp_fu_21465_p2[32'd13];

assign tmp_244_fu_3548_p3 = add_ln377_25_fu_3542_p2[32'd20];

assign tmp_245_fu_3562_p3 = add_ln1347_40_fu_3493_p2[32'd35];

assign tmp_246_fu_3588_p3 = add_ln1347_40_fu_3493_p2[32'd35];

assign tmp_247_fu_4307_p3 = select_ln346_106_fu_4300_p3[32'd20];

assign tmp_248_fu_4315_p3 = select_ln346_106_fu_4300_p3[32'd20];

assign tmp_249_fu_4357_p3 = select_ln346_108_fu_4349_p3[32'd20];

assign tmp_250_fu_4365_p3 = select_ln346_108_fu_4349_p3[32'd20];

assign tmp_251_fu_4407_p3 = select_ln346_110_fu_4399_p3[32'd20];

assign tmp_252_fu_4415_p3 = select_ln346_110_fu_4399_p3[32'd20];

assign tmp_253_fu_4457_p3 = select_ln346_112_fu_4449_p3[32'd20];

assign tmp_254_fu_4465_p3 = select_ln346_112_fu_4449_p3[32'd20];

assign tmp_255_fu_5820_p3 = add_ln1347_41_fu_5809_p2[32'd35];

assign tmp_256_fu_5838_p3 = add_ln810_19_fu_5815_p2[32'd34];

assign tmp_257_fu_5846_p3 = grp_fu_21530_p2[32'd13];

assign tmp_258_fu_5863_p3 = add_ln377_26_fu_5857_p2[32'd20];

assign tmp_259_fu_5877_p3 = add_ln1347_41_fu_5809_p2[32'd35];

assign tmp_260_fu_5903_p3 = add_ln1347_41_fu_5809_p2[32'd35];

assign tmp_261_fu_6501_p3 = add_ln1347_42_fu_6489_p2[32'd35];

assign tmp_262_fu_6519_p3 = add_ln810_20_fu_6495_p2[32'd34];

assign tmp_264_fu_6536_p3 = add_ln377_27_fu_6530_p2[32'd20];

assign tmp_265_fu_6556_p3 = add_ln1347_42_fu_6489_p2[32'd35];

assign tmp_266_fu_6582_p3 = add_ln1347_42_fu_6489_p2[32'd35];

assign tmp_267_fu_7122_p3 = select_ln346_118_fu_7116_p3[32'd20];

assign tmp_268_fu_7130_p3 = select_ln346_118_fu_7116_p3[32'd20];

assign tmp_269_fu_7172_p3 = select_ln346_120_fu_7164_p3[32'd20];

assign tmp_270_fu_7180_p3 = select_ln346_120_fu_7164_p3[32'd20];

assign tmp_271_fu_7239_p3 = add_ln1347_43_fu_7234_p2[32'd35];

assign tmp_272_fu_7257_p3 = add_ln1347_43_fu_7234_p2[32'd34];

assign tmp_273_fu_7265_p3 = grp_fu_21567_p2[32'd13];

assign tmp_274_fu_7282_p3 = add_ln377_28_fu_7276_p2[32'd20];

assign tmp_275_fu_7296_p3 = add_ln1347_43_fu_7234_p2[32'd35];

assign tmp_276_fu_7322_p3 = add_ln1347_43_fu_7234_p2[32'd35];

assign tmp_277_fu_7872_p3 = select_ln346_124_fu_7865_p3[32'd20];

assign tmp_278_fu_7880_p3 = select_ln346_124_fu_7865_p3[32'd20];

assign tmp_279_fu_7922_p3 = select_ln346_126_fu_7914_p3[32'd20];

assign tmp_280_fu_7930_p3 = select_ln346_126_fu_7914_p3[32'd20];

assign tmp_281_fu_7989_p3 = add_ln1347_44_fu_7984_p2[32'd35];

assign tmp_282_fu_8007_p3 = add_ln1347_44_fu_7984_p2[32'd34];

assign tmp_283_fu_8015_p3 = grp_fu_21582_p2[32'd13];

assign tmp_284_fu_8032_p3 = add_ln377_29_fu_8026_p2[32'd20];

assign tmp_285_fu_8046_p3 = add_ln1347_44_fu_7984_p2[32'd35];

assign tmp_286_fu_8072_p3 = add_ln1347_44_fu_7984_p2[32'd35];

assign tmp_287_fu_10286_p3 = sub_ln1348_fu_10281_p2[32'd21];

assign tmp_288_fu_10298_p3 = sub_ln1348_fu_10281_p2[32'd20];

assign tmp_289_fu_9564_p3 = sub_ln1348_18_fu_9559_p2[32'd21];

assign tmp_290_fu_9576_p3 = sub_ln1348_18_fu_9559_p2[32'd20];

assign tmp_291_fu_8663_p3 = sub_ln1348_19_fu_8658_p2[32'd21];

assign tmp_292_fu_8675_p3 = sub_ln1348_19_fu_8658_p2[32'd20];

assign tmp_293_fu_10366_p3 = grp_fu_21618_p2[32'd33];

assign tmp_294_fu_10386_p3 = grp_fu_21618_p2[32'd33];

assign tmp_295_fu_10393_p3 = grp_fu_21618_p2[32'd13];

assign tmp_296_fu_10410_p3 = add_ln377_30_fu_10404_p2[32'd20];

assign tmp_297_fu_10430_p3 = grp_fu_21618_p2[32'd33];

assign tmp_298_fu_10455_p3 = grp_fu_21618_p2[32'd33];

assign tmp_299_fu_10936_p3 = add_ln1347_45_fu_10924_p2[32'd35];

assign tmp_300_fu_10954_p3 = add_ln810_21_fu_10930_p2[32'd34];

assign tmp_302_fu_10971_p3 = add_ln377_31_fu_10965_p2[32'd20];

assign tmp_303_fu_10991_p3 = add_ln1347_45_fu_10924_p2[32'd35];

assign tmp_304_fu_11017_p3 = add_ln1347_45_fu_10924_p2[32'd35];

assign tmp_305_fu_11611_p3 = add_ln1347_46_fu_11599_p2[32'd35];

assign tmp_306_fu_11629_p3 = add_ln810_22_fu_11605_p2[32'd34];

assign tmp_308_fu_11646_p3 = add_ln377_32_fu_11640_p2[32'd20];

assign tmp_309_fu_11666_p3 = add_ln1347_46_fu_11599_p2[32'd35];

assign tmp_310_fu_11692_p3 = add_ln1347_46_fu_11599_p2[32'd35];

assign tmp_311_fu_10556_p3 = grp_fu_21630_p2[32'd30];

assign tmp_312_fu_10576_p3 = grp_fu_21630_p2[32'd30];

assign tmp_313_fu_10583_p3 = grp_fu_21630_p2[32'd13];

assign tmp_314_fu_10600_p3 = add_ln377_33_fu_10594_p2[32'd17];

assign tmp_315_fu_10620_p3 = grp_fu_21630_p2[32'd30];

assign tmp_316_fu_10645_p3 = grp_fu_21630_p2[32'd30];

assign tmp_317_fu_11166_p3 = add_ln1347_47_fu_11154_p2[32'd35];

assign tmp_318_fu_11184_p3 = add_ln810_23_fu_11160_p2[32'd34];

assign tmp_320_fu_11201_p3 = add_ln377_34_fu_11195_p2[32'd20];

assign tmp_321_fu_11221_p3 = add_ln1347_47_fu_11154_p2[32'd35];

assign tmp_322_fu_11247_p3 = add_ln1347_47_fu_11154_p2[32'd35];

assign tmp_323_fu_11807_p3 = add_ln1347_48_fu_11795_p2[32'd35];

assign tmp_324_fu_11825_p3 = add_ln810_24_fu_11801_p2[32'd34];

assign tmp_326_fu_11842_p3 = add_ln377_35_fu_11836_p2[32'd20];

assign tmp_327_fu_11862_p3 = add_ln1347_48_fu_11795_p2[32'd35];

assign tmp_328_fu_11888_p3 = add_ln1347_48_fu_11795_p2[32'd35];

assign tmp_329_fu_10730_p3 = grp_fu_21642_p2[32'd29];

assign tmp_330_fu_10750_p3 = grp_fu_21642_p2[32'd29];

assign tmp_331_fu_10757_p3 = grp_fu_21642_p2[32'd13];

assign tmp_332_fu_10774_p3 = add_ln377_36_fu_10768_p2[32'd16];

assign tmp_333_fu_10794_p3 = grp_fu_21642_p2[32'd29];

assign tmp_334_fu_10819_p3 = grp_fu_21642_p2[32'd29];

assign tmp_335_fu_11415_p3 = add_ln1347_49_fu_11403_p2[32'd35];

assign tmp_336_fu_11433_p3 = add_ln810_25_fu_11409_p2[32'd34];

assign tmp_338_fu_11450_p3 = add_ln377_37_fu_11444_p2[32'd20];

assign tmp_339_fu_11470_p3 = add_ln1347_49_fu_11403_p2[32'd35];

assign tmp_340_fu_11496_p3 = add_ln1347_49_fu_11403_p2[32'd35];

assign tmp_341_fu_12013_p3 = add_ln1347_50_fu_12002_p2[32'd35];

assign tmp_342_fu_12031_p3 = add_ln810_26_fu_12008_p2[32'd34];

assign tmp_344_fu_12048_p3 = add_ln377_38_fu_12042_p2[32'd20];

assign tmp_345_fu_12068_p3 = add_ln1347_50_fu_12002_p2[32'd35];

assign tmp_346_fu_12094_p3 = add_ln1347_50_fu_12002_p2[32'd35];

assign tmp_347_fu_13111_p3 = grp_fu_21654_p2[32'd34];

assign tmp_348_fu_13127_p3 = grp_fu_21654_p2[32'd34];

assign tmp_349_fu_13134_p3 = grp_fu_21654_p2[32'd13];

assign tmp_350_fu_13151_p3 = add_ln377_39_fu_13145_p2[32'd20];

assign tmp_351_fu_13171_p3 = grp_fu_21654_p2[32'd34];

assign tmp_352_fu_13196_p3 = grp_fu_21654_p2[32'd34];

assign tmp_353_fu_14944_p3 = select_ln346_153_fu_14938_p3[32'd20];

assign tmp_354_fu_14952_p3 = select_ln346_153_fu_14938_p3[32'd20];

assign tmp_355_fu_14994_p3 = select_ln346_155_fu_14986_p3[32'd20];

assign tmp_356_fu_15002_p3 = select_ln346_155_fu_14986_p3[32'd20];

assign tmp_357_fu_13281_p3 = grp_fu_21666_p2[32'd27];

assign tmp_358_fu_13301_p3 = grp_fu_21666_p2[32'd27];

assign tmp_359_fu_13308_p3 = grp_fu_21666_p2[32'd13];

assign tmp_360_fu_13325_p3 = add_ln377_40_fu_13319_p2[32'd14];

assign tmp_361_fu_13345_p3 = grp_fu_21666_p2[32'd27];

assign tmp_362_fu_13370_p3 = grp_fu_21666_p2[32'd27];

assign tmp_363_fu_15062_p3 = select_ln346_159_fu_15055_p3[32'd20];

assign tmp_364_fu_15070_p3 = select_ln346_159_fu_15055_p3[32'd20];

assign tmp_365_fu_15112_p3 = select_ln346_161_fu_15104_p3[32'd20];

assign tmp_366_fu_15120_p3 = select_ln346_161_fu_15104_p3[32'd20];

assign tmp_367_fu_13455_p3 = grp_fu_21678_p2[32'd34];

assign tmp_368_fu_13471_p3 = grp_fu_21678_p2[32'd34];

assign tmp_369_fu_13478_p3 = grp_fu_21678_p2[32'd13];

assign tmp_36_fu_1337_p3 = add_ln813_fu_1331_p2[32'd20];

assign tmp_370_fu_13495_p3 = add_ln377_41_fu_13489_p2[32'd20];

assign tmp_371_fu_13515_p3 = grp_fu_21678_p2[32'd34];

assign tmp_372_fu_13540_p3 = grp_fu_21678_p2[32'd34];

assign tmp_373_fu_15188_p3 = add_ln1347_51_fu_15177_p2[32'd35];

assign tmp_374_fu_15206_p3 = add_ln810_27_fu_15183_p2[32'd34];

assign tmp_375_fu_15214_p3 = grp_fu_21802_p2[32'd13];

assign tmp_376_fu_15231_p3 = add_ln377_42_fu_15225_p2[32'd20];

assign tmp_377_fu_15245_p3 = add_ln1347_51_fu_15177_p2[32'd35];

assign tmp_378_fu_15271_p3 = add_ln1347_51_fu_15177_p2[32'd35];

assign tmp_379_fu_17173_p3 = select_ln346_167_fu_17166_p3[32'd20];

assign tmp_37_fu_1393_p3 = add_ln1347_1_fu_1387_p2[32'd21];

assign tmp_380_fu_17181_p3 = select_ln346_167_fu_17166_p3[32'd20];

assign tmp_381_fu_13641_p3 = grp_fu_21690_p2[32'd28];

assign tmp_382_fu_13661_p3 = grp_fu_21690_p2[32'd28];

assign tmp_383_fu_13668_p3 = grp_fu_21690_p2[32'd13];

assign tmp_384_fu_13685_p3 = add_ln377_43_fu_13679_p2[32'd15];

assign tmp_385_fu_13705_p3 = grp_fu_21690_p2[32'd28];

assign tmp_386_fu_13730_p3 = grp_fu_21690_p2[32'd28];

assign tmp_387_fu_15380_p3 = add_ln1347_52_fu_15368_p2[32'd35];

assign tmp_388_fu_15398_p3 = add_ln810_28_fu_15374_p2[32'd34];

assign tmp_389_fu_15406_p3 = grp_fu_21810_p2[32'd13];

assign tmp_38_fu_1407_p3 = add_ln813_1_fu_1401_p2[32'd20];

assign tmp_390_fu_15423_p3 = add_ln377_44_fu_15417_p2[32'd20];

assign tmp_391_fu_15437_p3 = add_ln1347_52_fu_15368_p2[32'd35];

assign tmp_392_fu_15463_p3 = add_ln1347_52_fu_15368_p2[32'd35];

assign tmp_393_fu_17261_p3 = select_ln346_173_fu_17254_p3[32'd20];

assign tmp_394_fu_17269_p3 = select_ln346_173_fu_17254_p3[32'd20];

assign tmp_395_fu_13815_p3 = grp_fu_21702_p2[32'd33];

assign tmp_396_fu_13835_p3 = grp_fu_21702_p2[32'd33];

assign tmp_397_fu_13842_p3 = grp_fu_21702_p2[32'd13];

assign tmp_398_fu_13859_p3 = add_ln377_45_fu_13853_p2[32'd20];

assign tmp_399_fu_13879_p3 = grp_fu_21702_p2[32'd33];

assign tmp_39_fu_1471_p3 = add_ln1347_2_fu_1465_p2[32'd21];

assign tmp_400_fu_13904_p3 = grp_fu_21702_p2[32'd33];

assign tmp_401_fu_15550_p3 = add_ln1347_53_fu_15539_p2[32'd35];

assign tmp_402_fu_15568_p3 = add_ln810_29_fu_15545_p2[32'd34];

assign tmp_404_fu_15585_p3 = add_ln377_46_fu_15579_p2[32'd20];

assign tmp_405_fu_15605_p3 = add_ln1347_53_fu_15539_p2[32'd35];

assign tmp_406_fu_15631_p3 = add_ln1347_53_fu_15539_p2[32'd35];

assign tmp_407_fu_17336_p3 = add_ln1347_54_fu_17325_p2[32'd35];

assign tmp_408_fu_17354_p3 = add_ln810_30_fu_17331_p2[32'd34];

assign tmp_40_fu_1485_p3 = add_ln813_2_fu_1479_p2[32'd20];

assign tmp_410_fu_17371_p3 = add_ln377_47_fu_17365_p2[32'd20];

assign tmp_411_fu_17391_p3 = add_ln1347_54_fu_17325_p2[32'd35];

assign tmp_412_fu_17417_p3 = add_ln1347_54_fu_17325_p2[32'd35];

assign tmp_413_fu_14012_p3 = grp_fu_21721_p2[32'd29];

assign tmp_414_fu_14032_p3 = grp_fu_21721_p2[32'd29];

assign tmp_415_fu_14039_p3 = grp_fu_21721_p2[32'd13];

assign tmp_416_fu_14056_p3 = add_ln377_48_fu_14050_p2[32'd16];

assign tmp_417_fu_14076_p3 = grp_fu_21721_p2[32'd29];

assign tmp_418_fu_14101_p3 = grp_fu_21721_p2[32'd29];

assign tmp_419_fu_15787_p3 = add_ln1347_55_fu_15775_p2[32'd35];

assign tmp_41_fu_1623_p3 = add_ln1347_3_fu_1617_p2[32'd21];

assign tmp_420_fu_15805_p3 = add_ln810_31_fu_15781_p2[32'd34];

assign tmp_422_fu_15822_p3 = add_ln377_49_fu_15816_p2[32'd20];

assign tmp_423_fu_15842_p3 = add_ln1347_55_fu_15775_p2[32'd35];

assign tmp_424_fu_15868_p3 = add_ln1347_55_fu_15775_p2[32'd35];

assign tmp_425_fu_17548_p3 = add_ln1347_56_fu_17536_p2[32'd35];

assign tmp_426_fu_17566_p3 = add_ln810_32_fu_17542_p2[32'd34];

assign tmp_428_fu_17583_p3 = add_ln377_50_fu_17577_p2[32'd20];

assign tmp_429_fu_17603_p3 = add_ln1347_56_fu_17536_p2[32'd35];

assign tmp_42_fu_1637_p3 = add_ln813_3_fu_1631_p2[32'd20];

assign tmp_430_fu_17629_p3 = add_ln1347_56_fu_17536_p2[32'd35];

assign tmp_431_fu_15977_p3 = grp_fu_21833_p2[32'd34];

assign tmp_432_fu_15993_p3 = grp_fu_21833_p2[32'd34];

assign tmp_433_fu_16000_p3 = grp_fu_21833_p2[32'd13];

assign tmp_434_fu_16017_p3 = add_ln377_51_fu_16011_p2[32'd20];

assign tmp_435_fu_16037_p3 = grp_fu_21833_p2[32'd34];

assign tmp_436_fu_16062_p3 = grp_fu_21833_p2[32'd34];

assign tmp_437_fu_17744_p3 = select_ln346_189_fu_17738_p3[32'd20];

assign tmp_438_fu_17752_p3 = select_ln346_189_fu_17738_p3[32'd20];

assign tmp_439_fu_17794_p3 = select_ln346_191_fu_17786_p3[32'd20];

assign tmp_43_fu_1541_p3 = add_ln1347_4_fu_1535_p2[32'd21];

assign tmp_440_fu_17802_p3 = select_ln346_191_fu_17786_p3[32'd20];

assign tmp_441_fu_16147_p3 = grp_fu_21844_p2[32'd27];

assign tmp_442_fu_16167_p3 = grp_fu_21844_p2[32'd27];

assign tmp_443_fu_16174_p3 = grp_fu_21844_p2[32'd13];

assign tmp_444_fu_16191_p3 = add_ln377_52_fu_16185_p2[32'd14];

assign tmp_445_fu_16211_p3 = grp_fu_21844_p2[32'd27];

assign tmp_446_fu_16236_p3 = grp_fu_21844_p2[32'd27];

assign tmp_447_fu_17862_p3 = select_ln346_195_fu_17855_p3[32'd20];

assign tmp_448_fu_17870_p3 = select_ln346_195_fu_17855_p3[32'd20];

assign tmp_449_fu_17912_p3 = select_ln346_197_fu_17904_p3[32'd20];

assign tmp_44_fu_1555_p3 = add_ln813_4_fu_1549_p2[32'd20];

assign tmp_450_fu_17920_p3 = select_ln346_197_fu_17904_p3[32'd20];

assign tmp_451_fu_14193_p3 = grp_fu_21740_p2[32'd34];

assign tmp_452_fu_14209_p3 = grp_fu_21740_p2[32'd34];

assign tmp_453_fu_14216_p3 = grp_fu_21740_p2[32'd13];

assign tmp_454_fu_14233_p3 = add_ln377_53_fu_14227_p2[32'd20];

assign tmp_455_fu_14253_p3 = grp_fu_21740_p2[32'd34];

assign tmp_456_fu_14278_p3 = grp_fu_21740_p2[32'd34];

assign tmp_457_fu_16346_p3 = add_ln1347_57_fu_16335_p2[32'd35];

assign tmp_458_fu_16364_p3 = add_ln810_33_fu_16341_p2[32'd34];

assign tmp_459_fu_16372_p3 = grp_fu_21855_p2[32'd13];

assign tmp_45_fu_1693_p3 = add_ln1347_5_fu_1687_p2[32'd21];

assign tmp_460_fu_16389_p3 = add_ln377_54_fu_16383_p2[32'd20];

assign tmp_461_fu_16403_p3 = add_ln1347_57_fu_16335_p2[32'd35];

assign tmp_462_fu_16429_p3 = add_ln1347_57_fu_16335_p2[32'd35];

assign tmp_463_fu_18001_p3 = select_ln346_203_fu_17994_p3[32'd20];

assign tmp_464_fu_18009_p3 = select_ln346_203_fu_17994_p3[32'd20];

assign tmp_465_fu_14379_p3 = grp_fu_21752_p2[32'd28];

assign tmp_466_fu_14399_p3 = grp_fu_21752_p2[32'd28];

assign tmp_467_fu_14406_p3 = grp_fu_21752_p2[32'd13];

assign tmp_468_fu_14423_p3 = add_ln377_55_fu_14417_p2[32'd15];

assign tmp_469_fu_14443_p3 = grp_fu_21752_p2[32'd28];

assign tmp_46_fu_1707_p3 = add_ln813_5_fu_1701_p2[32'd20];

assign tmp_470_fu_14468_p3 = grp_fu_21752_p2[32'd28];

assign tmp_471_fu_16538_p3 = add_ln1347_58_fu_16526_p2[32'd35];

assign tmp_472_fu_16556_p3 = add_ln810_34_fu_16532_p2[32'd34];

assign tmp_473_fu_16564_p3 = grp_fu_21863_p2[32'd13];

assign tmp_474_fu_16581_p3 = add_ln377_56_fu_16575_p2[32'd20];

assign tmp_475_fu_16595_p3 = add_ln1347_58_fu_16526_p2[32'd35];

assign tmp_476_fu_16621_p3 = add_ln1347_58_fu_16526_p2[32'd35];

assign tmp_477_fu_18089_p3 = select_ln346_209_fu_18082_p3[32'd20];

assign tmp_478_fu_18097_p3 = select_ln346_209_fu_18082_p3[32'd20];

assign tmp_479_fu_14553_p3 = grp_fu_21764_p2[32'd33];

assign tmp_47_fu_1851_p3 = add_ln1347_6_fu_1845_p2[32'd21];

assign tmp_480_fu_14573_p3 = grp_fu_21764_p2[32'd33];

assign tmp_481_fu_14580_p3 = grp_fu_21764_p2[32'd13];

assign tmp_482_fu_14597_p3 = add_ln377_57_fu_14591_p2[32'd20];

assign tmp_483_fu_14617_p3 = grp_fu_21764_p2[32'd33];

assign tmp_484_fu_14642_p3 = grp_fu_21764_p2[32'd33];

assign tmp_485_fu_16708_p3 = add_ln1347_59_fu_16697_p2[32'd35];

assign tmp_486_fu_16726_p3 = add_ln810_35_fu_16703_p2[32'd34];

assign tmp_488_fu_16743_p3 = add_ln377_58_fu_16737_p2[32'd20];

assign tmp_489_fu_16763_p3 = add_ln1347_59_fu_16697_p2[32'd35];

assign tmp_48_fu_1865_p3 = add_ln813_6_fu_1859_p2[32'd20];

assign tmp_490_fu_16789_p3 = add_ln1347_59_fu_16697_p2[32'd35];

assign tmp_491_fu_18164_p3 = add_ln1347_60_fu_18153_p2[32'd35];

assign tmp_492_fu_18182_p3 = add_ln810_36_fu_18159_p2[32'd34];

assign tmp_494_fu_18199_p3 = add_ln377_59_fu_18193_p2[32'd20];

assign tmp_495_fu_18219_p3 = add_ln1347_60_fu_18153_p2[32'd35];

assign tmp_496_fu_18245_p3 = add_ln1347_60_fu_18153_p2[32'd35];

assign tmp_497_fu_14750_p3 = grp_fu_21783_p2[32'd29];

assign tmp_498_fu_14770_p3 = grp_fu_21783_p2[32'd29];

assign tmp_499_fu_14777_p3 = grp_fu_21783_p2[32'd13];

assign tmp_49_fu_1921_p3 = add_ln1347_7_fu_1915_p2[32'd21];

assign tmp_500_fu_14794_p3 = add_ln377_60_fu_14788_p2[32'd16];

assign tmp_501_fu_14814_p3 = grp_fu_21783_p2[32'd29];

assign tmp_502_fu_14839_p3 = grp_fu_21783_p2[32'd29];

assign tmp_503_fu_16945_p3 = add_ln1347_61_fu_16933_p2[32'd35];

assign tmp_504_fu_16963_p3 = add_ln810_37_fu_16939_p2[32'd34];

assign tmp_506_fu_16980_p3 = add_ln377_61_fu_16974_p2[32'd20];

assign tmp_507_fu_17000_p3 = add_ln1347_61_fu_16933_p2[32'd35];

assign tmp_508_fu_17026_p3 = add_ln1347_61_fu_16933_p2[32'd35];

assign tmp_509_fu_18376_p3 = add_ln1347_62_fu_18364_p2[32'd35];

assign tmp_50_fu_1935_p3 = add_ln813_7_fu_1929_p2[32'd20];

assign tmp_510_fu_18394_p3 = add_ln810_38_fu_18370_p2[32'd34];

assign tmp_512_fu_18411_p3 = add_ln377_62_fu_18405_p2[32'd20];

assign tmp_513_fu_18431_p3 = add_ln1347_62_fu_18364_p2[32'd35];

assign tmp_514_fu_18457_p3 = add_ln1347_62_fu_18364_p2[32'd35];

assign tmp_515_fu_12240_p3 = select_ln346_139_fu_12187_p3[32'd20];

assign tmp_516_fu_12248_p3 = select_ln346_139_fu_12187_p3[32'd20];

assign tmp_517_fu_12290_p3 = select_ln346_225_fu_12282_p3[32'd20];

assign tmp_518_fu_12298_p3 = select_ln346_225_fu_12282_p3[32'd20];

assign tmp_519_fu_12340_p3 = select_ln346_227_fu_12332_p3[32'd20];

assign tmp_51_fu_2192_p3 = add_ln1347_8_fu_2186_p2[32'd21];

assign tmp_520_fu_12348_p3 = select_ln346_227_fu_12332_p3[32'd20];

assign tmp_521_fu_12391_p3 = select_ln346_145_fu_12206_p3[32'd20];

assign tmp_522_fu_12399_p3 = select_ln346_145_fu_12206_p3[32'd20];

assign tmp_523_fu_12407_p3 = select_ln346_145_fu_12206_p3[32'd20];

assign tmp_524_fu_12473_p3 = select_ln346_231_fu_12465_p3[32'd20];

assign tmp_525_fu_12481_p3 = select_ln346_231_fu_12465_p3[32'd20];

assign tmp_526_fu_12548_p3 = select_ln346_151_fu_12531_p3[32'd20];

assign tmp_527_fu_12556_p3 = select_ln346_151_fu_12531_p3[32'd20];

assign tmp_528_fu_12564_p3 = select_ln346_151_fu_12531_p3[32'd20];

assign tmp_529_fu_12648_p3 = sub_ln1273_6_fu_12642_p2[32'd35];

assign tmp_52_fu_2206_p3 = add_ln813_8_fu_2200_p2[32'd20];

assign tmp_530_fu_12666_p3 = sub_ln1273_6_fu_12642_p2[32'd34];

assign tmp_531_fu_12674_p3 = sub_ln1273_6_fu_12642_p2[32'd35];

assign tmp_532_fu_12740_p3 = select_ln346_237_fu_12732_p3[32'd20];

assign tmp_533_fu_12748_p3 = select_ln346_237_fu_12732_p3[32'd20];

assign tmp_534_fu_12790_p3 = select_ln346_239_fu_12782_p3[32'd20];

assign tmp_535_fu_12798_p3 = select_ln346_239_fu_12782_p3[32'd20];

assign tmp_536_fu_12869_p3 = sub_ln1273_7_fu_12863_p2[32'd35];

assign tmp_537_fu_12887_p3 = sub_ln1273_7_fu_12863_p2[32'd34];

assign tmp_538_fu_12895_p3 = sub_ln1273_7_fu_12863_p2[32'd35];

assign tmp_539_fu_12961_p3 = select_ln346_243_fu_12953_p3[32'd20];

assign tmp_53_fu_2262_p3 = add_ln1347_9_fu_2256_p2[32'd21];

assign tmp_540_fu_12969_p3 = select_ln346_243_fu_12953_p3[32'd20];

assign tmp_541_fu_13018_p3 = sub_ln1273_8_fu_13012_p2[32'd35];

assign tmp_542_fu_13036_p3 = sub_ln1273_8_fu_13012_p2[32'd34];

assign tmp_543_fu_13044_p3 = sub_ln1273_8_fu_13012_p2[32'd35];

assign tmp_544_fu_18573_p3 = add_ln1347_63_fu_18567_p2[32'd21];

assign tmp_545_fu_18587_p3 = add_ln813_18_fu_18581_p2[32'd20];

assign tmp_546_fu_18644_p3 = add_ln1347_64_fu_18638_p2[32'd21];

assign tmp_547_fu_18658_p3 = add_ln813_19_fu_18652_p2[32'd20];

assign tmp_548_fu_18749_p3 = add_ln1347_65_fu_18743_p2[32'd21];

assign tmp_549_fu_18763_p3 = add_ln813_20_fu_18757_p2[32'd20];

assign tmp_54_fu_2276_p3 = add_ln813_9_fu_2270_p2[32'd20];

assign tmp_550_fu_18820_p3 = add_ln1347_66_fu_18814_p2[32'd21];

assign tmp_551_fu_18834_p3 = add_ln813_21_fu_18828_p2[32'd20];

assign tmp_552_fu_18925_p3 = add_ln1347_67_fu_18919_p2[32'd21];

assign tmp_553_fu_18939_p3 = add_ln813_22_fu_18933_p2[32'd20];

assign tmp_554_fu_18996_p3 = add_ln1347_68_fu_18990_p2[32'd21];

assign tmp_555_fu_19010_p3 = add_ln813_23_fu_19004_p2[32'd20];

assign tmp_556_fu_19101_p3 = add_ln1347_69_fu_19095_p2[32'd21];

assign tmp_557_fu_19115_p3 = add_ln813_24_fu_19109_p2[32'd20];

assign tmp_558_fu_19172_p3 = add_ln1347_70_fu_19166_p2[32'd21];

assign tmp_559_fu_19186_p3 = add_ln813_25_fu_19180_p2[32'd20];

assign tmp_55_fu_2945_p3 = add_ln1347_10_fu_2939_p2[32'd21];

assign tmp_560_fu_19277_p3 = add_ln1347_71_fu_19271_p2[32'd21];

assign tmp_561_fu_19291_p3 = add_ln813_26_fu_19285_p2[32'd20];

assign tmp_562_fu_19348_p3 = add_ln1347_72_fu_19342_p2[32'd21];

assign tmp_563_fu_19362_p3 = add_ln813_27_fu_19356_p2[32'd20];

assign tmp_564_fu_19453_p3 = add_ln1347_73_fu_19447_p2[32'd21];

assign tmp_565_fu_19467_p3 = add_ln813_28_fu_19461_p2[32'd20];

assign tmp_566_fu_19524_p3 = add_ln1347_74_fu_19518_p2[32'd21];

assign tmp_567_fu_19538_p3 = add_ln813_29_fu_19532_p2[32'd20];

assign tmp_568_fu_19629_p3 = add_ln1347_75_fu_19623_p2[32'd21];

assign tmp_569_fu_19643_p3 = add_ln813_30_fu_19637_p2[32'd20];

assign tmp_56_fu_2959_p3 = add_ln813_10_fu_2953_p2[32'd20];

assign tmp_570_fu_19700_p3 = add_ln1347_76_fu_19694_p2[32'd21];

assign tmp_571_fu_19714_p3 = add_ln813_31_fu_19708_p2[32'd20];

assign tmp_572_fu_19805_p3 = add_ln1347_77_fu_19799_p2[32'd21];

assign tmp_573_fu_19819_p3 = add_ln813_32_fu_19813_p2[32'd20];

assign tmp_574_fu_19876_p3 = add_ln1347_78_fu_19870_p2[32'd21];

assign tmp_575_fu_19890_p3 = add_ln813_33_fu_19884_p2[32'd20];

assign tmp_576_fu_19981_p3 = add_ln1347_79_fu_19975_p2[32'd21];

assign tmp_577_fu_19995_p3 = add_ln813_34_fu_19989_p2[32'd20];

assign tmp_578_fu_20052_p3 = add_ln1347_80_fu_20046_p2[32'd21];

assign tmp_579_fu_20066_p3 = add_ln813_35_fu_20060_p2[32'd20];

assign tmp_57_fu_3015_p3 = add_ln1347_11_fu_3009_p2[32'd21];

assign tmp_580_fu_20156_p3 = add_ln1347_81_fu_20150_p2[32'd21];

assign tmp_581_fu_20169_p3 = add_ln813_36_fu_20164_p2[32'd20];

assign tmp_582_fu_20225_p3 = add_ln1347_82_fu_20219_p2[32'd21];

assign tmp_583_fu_20238_p3 = add_ln813_37_fu_20233_p2[32'd20];

assign tmp_584_fu_20294_p3 = add_ln1347_83_fu_20288_p2[32'd21];

assign tmp_585_fu_20307_p3 = add_ln813_38_fu_20302_p2[32'd20];

assign tmp_586_fu_20363_p3 = add_ln1347_84_fu_20357_p2[32'd21];

assign tmp_587_fu_20376_p3 = add_ln813_39_fu_20371_p2[32'd20];

assign tmp_588_fu_20432_p3 = add_ln1347_85_fu_20426_p2[32'd21];

assign tmp_589_fu_20445_p3 = add_ln813_40_fu_20440_p2[32'd20];

assign tmp_58_fu_3029_p3 = add_ln813_11_fu_3023_p2[32'd20];

assign tmp_590_fu_20501_p3 = add_ln1347_86_fu_20495_p2[32'd21];

assign tmp_591_fu_20514_p3 = add_ln813_41_fu_20509_p2[32'd20];

assign tmp_592_fu_20570_p3 = add_ln1347_87_fu_20564_p2[32'd21];

assign tmp_593_fu_20583_p3 = add_ln813_42_fu_20578_p2[32'd20];

assign tmp_594_fu_20639_p3 = add_ln1347_88_fu_20633_p2[32'd21];

assign tmp_595_fu_20652_p3 = add_ln813_43_fu_20647_p2[32'd20];

assign tmp_596_fu_20708_p3 = add_ln1347_89_fu_20702_p2[32'd21];

assign tmp_597_fu_20721_p3 = add_ln813_44_fu_20716_p2[32'd20];

assign tmp_598_fu_20777_p3 = add_ln1347_90_fu_20771_p2[32'd21];

assign tmp_599_fu_20790_p3 = add_ln813_45_fu_20785_p2[32'd20];

assign tmp_59_fu_3664_p3 = add_ln1347_12_fu_3658_p2[32'd21];

assign tmp_600_fu_20846_p3 = add_ln1347_91_fu_20840_p2[32'd21];

assign tmp_601_fu_20859_p3 = add_ln813_46_fu_20854_p2[32'd20];

assign tmp_602_fu_20915_p3 = add_ln1347_92_fu_20909_p2[32'd21];

assign tmp_603_fu_20928_p3 = add_ln813_47_fu_20923_p2[32'd20];

assign tmp_604_fu_20984_p3 = add_ln1347_93_fu_20978_p2[32'd21];

assign tmp_605_fu_20997_p3 = add_ln813_48_fu_20992_p2[32'd20];

assign tmp_606_fu_21053_p3 = add_ln1347_94_fu_21047_p2[32'd21];

assign tmp_607_fu_21066_p3 = add_ln813_49_fu_21061_p2[32'd20];

assign tmp_608_fu_21122_p3 = add_ln1347_95_fu_21116_p2[32'd21];

assign tmp_609_fu_21135_p3 = add_ln813_50_fu_21130_p2[32'd20];

assign tmp_60_fu_3678_p3 = add_ln813_12_fu_3672_p2[32'd20];

assign tmp_610_fu_21191_p3 = add_ln1347_96_fu_21185_p2[32'd21];

assign tmp_611_fu_21204_p3 = add_ln813_51_fu_21199_p2[32'd20];

assign tmp_612_fu_21260_p3 = add_ln1347_97_fu_21254_p2[32'd21];

assign tmp_613_fu_21273_p3 = add_ln813_52_fu_21268_p2[32'd20];

assign tmp_614_fu_21329_p3 = add_ln1347_98_fu_21323_p2[32'd21];

assign tmp_615_fu_21342_p3 = add_ln813_53_fu_21337_p2[32'd20];

assign tmp_61_fu_3734_p3 = add_ln1347_13_fu_3728_p2[32'd21];

assign tmp_62_fu_3748_p3 = add_ln813_13_fu_3742_p2[32'd20];

assign tmp_63_fu_4521_p3 = add_ln1347_14_fu_4515_p2[32'd21];

assign tmp_64_fu_4535_p3 = add_ln813_14_fu_4529_p2[32'd20];

assign tmp_65_fu_4591_p3 = add_ln1347_15_fu_4585_p2[32'd21];

assign tmp_66_fu_4605_p3 = add_ln813_15_fu_4599_p2[32'd20];

assign tmp_67_fu_5156_p3 = add_ln1347_16_fu_5150_p2[32'd21];

assign tmp_68_fu_5170_p3 = add_ln813_16_fu_5164_p2[32'd20];

assign tmp_69_fu_5226_p3 = add_ln1347_17_fu_5220_p2[32'd21];

assign tmp_70_fu_5240_p3 = add_ln813_17_fu_5234_p2[32'd20];

assign tmp_71_fu_1977_p3 = grp_fu_21385_p2[32'd34];

assign tmp_72_fu_1993_p3 = grp_fu_21385_p2[32'd34];

assign tmp_73_fu_2000_p3 = grp_fu_21385_p2[32'd13];

assign tmp_74_fu_2017_p3 = add_ln377_fu_2011_p2[32'd20];

assign tmp_75_fu_2037_p3 = grp_fu_21385_p2[32'd34];

assign tmp_76_fu_2062_p3 = grp_fu_21385_p2[32'd34];

assign tmp_77_fu_2347_p3 = add_ln1347_18_fu_2335_p2[32'd35];

assign tmp_78_fu_2365_p3 = add_ln810_fu_2341_p2[32'd34];

assign tmp_80_fu_2382_p3 = add_ln377_1_fu_2376_p2[32'd20];

assign tmp_81_fu_2402_p3 = add_ln1347_18_fu_2335_p2[32'd35];

assign tmp_82_fu_2428_p3 = add_ln1347_18_fu_2335_p2[32'd35];

assign tmp_83_fu_3096_p3 = add_ln1347_19_fu_3085_p2[32'd35];

assign tmp_84_fu_3114_p3 = add_ln810_1_fu_3091_p2[32'd34];

assign tmp_86_fu_3131_p3 = add_ln377_2_fu_3125_p2[32'd20];

assign tmp_87_fu_3151_p3 = add_ln1347_19_fu_3085_p2[32'd35];

assign tmp_88_fu_3177_p3 = add_ln1347_19_fu_3085_p2[32'd35];

assign tmp_89_fu_3849_p3 = add_ln1347_20_fu_3837_p2[32'd35];

assign tmp_90_fu_3867_p3 = add_ln810_2_fu_3843_p2[32'd34];

assign tmp_92_fu_3884_p3 = add_ln377_3_fu_3878_p2[32'd20];

assign tmp_93_fu_3904_p3 = add_ln1347_20_fu_3837_p2[32'd35];

assign tmp_94_fu_3930_p3 = add_ln1347_20_fu_3837_p2[32'd35];

assign tmp_95_fu_4690_p3 = add_ln1347_21_fu_4678_p2[32'd35];

assign tmp_96_fu_4708_p3 = add_ln810_3_fu_4684_p2[32'd34];

assign tmp_98_fu_4725_p3 = add_ln377_4_fu_4719_p2[32'd20];

assign tmp_99_fu_4745_p3 = add_ln1347_21_fu_4678_p2[32'd35];

assign tmp_fu_1323_p3 = add_ln1347_fu_1317_p2[32'd21];

assign trunc_ln1273_10_fu_8749_p1 = select_ln302_23_fu_8709_p3[13:0];

assign trunc_ln1273_11_fu_9626_p1 = select_ln302_22_fu_9610_p3[5:0];

assign trunc_ln1273_12_fu_9638_p1 = select_ln302_22_fu_9610_p3[13:0];

assign trunc_ln1273_1_fu_1769_p3 = {{trunc_ln1273_6_fu_1765_p1}, {5'd0}};

assign trunc_ln1273_2_fu_1803_p3 = {{trunc_ln1273_7_fu_1799_p1}, {7'd0}};

assign trunc_ln1273_3_fu_1815_p3 = {{trunc_ln1273_8_fu_1811_p1}, {5'd0}};

assign trunc_ln1273_4_fu_8741_p3 = {{trunc_ln1273_9_fu_8737_p1}, {8'd0}};

assign trunc_ln1273_5_fu_9630_p3 = {{trunc_ln1273_11_fu_9626_p1}, {8'd0}};

assign trunc_ln1273_6_fu_1765_p1 = select_ln302_3_fu_1671_p3[8:0];

assign trunc_ln1273_7_fu_1799_p1 = select_ln302_5_fu_1741_p3[6:0];

assign trunc_ln1273_8_fu_1811_p1 = select_ln302_5_fu_1741_p3[8:0];

assign trunc_ln1273_9_fu_8737_p1 = select_ln302_23_fu_8709_p3[5:0];

assign trunc_ln1273_fu_1753_p1 = select_ln302_3_fu_1671_p3[6:0];

assign trunc_ln1649_10_fu_19581_p1 = temp5_q1[19:0];

assign trunc_ln1649_11_fu_19598_p1 = temp5_q0[19:0];

assign trunc_ln1649_12_fu_19757_p1 = temp5_q1[19:0];

assign trunc_ln1649_13_fu_19774_p1 = temp5_q0[19:0];

assign trunc_ln1649_14_fu_19933_p1 = temp5_q1[19:0];

assign trunc_ln1649_15_fu_19950_p1 = temp5_q0[19:0];

assign trunc_ln1649_16_fu_20109_p1 = temp5_q1[19:0];

assign trunc_ln1649_17_fu_20126_p1 = temp5_q0[19:0];

assign trunc_ln1649_1_fu_18718_p1 = temp5_q0[19:0];

assign trunc_ln1649_2_fu_18877_p1 = temp5_q1[19:0];

assign trunc_ln1649_3_fu_18894_p1 = temp5_q0[19:0];

assign trunc_ln1649_4_fu_19053_p1 = temp5_q1[19:0];

assign trunc_ln1649_5_fu_19070_p1 = temp5_q0[19:0];

assign trunc_ln1649_6_fu_19229_p1 = temp5_q1[19:0];

assign trunc_ln1649_7_fu_19246_p1 = temp5_q0[19:0];

assign trunc_ln1649_8_fu_19405_p1 = temp5_q1[19:0];

assign trunc_ln1649_9_fu_19422_p1 = temp5_q0[19:0];

assign trunc_ln1649_fu_18701_p1 = temp5_q1[19:0];

assign trunc_ln2_fu_1757_p3 = {{trunc_ln1273_fu_1753_p1}, {7'd0}};

assign trunc_ln813_18_fu_9572_p1 = sub_ln1348_18_fu_9559_p2[20:0];

assign trunc_ln813_19_fu_8671_p1 = sub_ln1348_19_fu_8658_p2[20:0];

assign trunc_ln813_fu_10294_p1 = sub_ln1348_fu_10281_p2[20:0];

assign trunc_ln818_10_fu_9333_p4 = {{add_ln810_10_fu_9319_p2[34:14]}};

assign trunc_ln818_11_fu_9694_p4 = {{add_ln1347_29_fu_9681_p2[34:14]}};

assign trunc_ln818_12_fu_10005_p4 = {{add_ln1347_30_fu_9992_p2[34:14]}};

assign trunc_ln818_13_fu_2559_p4 = {{grp_fu_21418_p2[34:14]}};

assign trunc_ln818_14_fu_3339_p4 = {{add_ln810_11_fu_3325_p2[34:14]}};

assign trunc_ln818_15_fu_4106_p4 = {{add_ln810_12_fu_4093_p2[34:14]}};

assign trunc_ln818_16_fu_4965_p4 = {{add_ln810_13_fu_4951_p2[34:14]}};

assign trunc_ln818_17_fu_5655_p4 = {{add_ln810_14_fu_5642_p2[34:14]}};

assign trunc_ln818_18_fu_6267_p4 = {{add_ln810_15_fu_6253_p2[34:14]}};

assign trunc_ln818_19_fu_6934_p4 = {{add_ln810_16_fu_6921_p2[34:14]}};

assign trunc_ln818_1_fu_2355_p4 = {{add_ln810_fu_2341_p2[34:14]}};

assign trunc_ln818_20_fu_7659_p4 = {{add_ln810_17_fu_7645_p2[34:14]}};

assign trunc_ln818_21_fu_8457_p4 = {{add_ln1347_38_fu_8444_p2[34:14]}};

assign trunc_ln818_22_fu_9137_p4 = {{add_ln1347_39_fu_9124_p2[34:14]}};

assign trunc_ln818_23_fu_2752_p4 = {{grp_fu_21437_p2[34:14]}};

assign trunc_ln818_24_fu_3513_p4 = {{add_ln810_18_fu_3499_p2[34:14]}};

assign trunc_ln818_25_fu_5828_p4 = {{add_ln810_19_fu_5815_p2[34:14]}};

assign trunc_ln818_26_fu_6509_p4 = {{add_ln810_20_fu_6495_p2[34:14]}};

assign trunc_ln818_27_fu_7247_p4 = {{add_ln1347_43_fu_7234_p2[34:14]}};

assign trunc_ln818_28_fu_7997_p4 = {{add_ln1347_44_fu_7984_p2[34:14]}};

assign trunc_ln818_29_fu_10373_p4 = {{grp_fu_21618_p2[33:14]}};

assign trunc_ln818_2_fu_3104_p4 = {{add_ln810_1_fu_3091_p2[34:14]}};

assign trunc_ln818_30_fu_10944_p4 = {{add_ln810_21_fu_10930_p2[34:14]}};

assign trunc_ln818_31_fu_11619_p4 = {{add_ln810_22_fu_11605_p2[34:14]}};

assign trunc_ln818_32_fu_10563_p4 = {{grp_fu_21630_p2[30:14]}};

assign trunc_ln818_33_fu_11174_p4 = {{add_ln810_23_fu_11160_p2[34:14]}};

assign trunc_ln818_34_fu_11815_p4 = {{add_ln810_24_fu_11801_p2[34:14]}};

assign trunc_ln818_35_fu_10737_p4 = {{grp_fu_21642_p2[29:14]}};

assign trunc_ln818_36_fu_11423_p4 = {{add_ln810_25_fu_11409_p2[34:14]}};

assign trunc_ln818_37_fu_12021_p4 = {{add_ln810_26_fu_12008_p2[34:14]}};

assign trunc_ln818_38_fu_13118_p4 = {{grp_fu_21654_p2[34:14]}};

assign trunc_ln818_39_fu_13288_p4 = {{grp_fu_21666_p2[27:14]}};

assign trunc_ln818_3_fu_3857_p4 = {{add_ln810_2_fu_3843_p2[34:14]}};

assign trunc_ln818_40_fu_13462_p4 = {{grp_fu_21678_p2[34:14]}};

assign trunc_ln818_41_fu_15196_p4 = {{add_ln810_27_fu_15183_p2[34:14]}};

assign trunc_ln818_42_fu_13648_p4 = {{grp_fu_21690_p2[28:14]}};

assign trunc_ln818_43_fu_15388_p4 = {{add_ln810_28_fu_15374_p2[34:14]}};

assign trunc_ln818_44_fu_13822_p4 = {{grp_fu_21702_p2[33:14]}};

assign trunc_ln818_45_fu_15558_p4 = {{add_ln810_29_fu_15545_p2[34:14]}};

assign trunc_ln818_46_fu_17344_p4 = {{add_ln810_30_fu_17331_p2[34:14]}};

assign trunc_ln818_47_fu_14019_p4 = {{grp_fu_21721_p2[29:14]}};

assign trunc_ln818_48_fu_15795_p4 = {{add_ln810_31_fu_15781_p2[34:14]}};

assign trunc_ln818_49_fu_17556_p4 = {{add_ln810_32_fu_17542_p2[34:14]}};

assign trunc_ln818_4_fu_4698_p4 = {{add_ln810_3_fu_4684_p2[34:14]}};

assign trunc_ln818_50_fu_15984_p4 = {{grp_fu_21833_p2[34:14]}};

assign trunc_ln818_51_fu_16154_p4 = {{grp_fu_21844_p2[27:14]}};

assign trunc_ln818_52_fu_14200_p4 = {{grp_fu_21740_p2[34:14]}};

assign trunc_ln818_53_fu_16354_p4 = {{add_ln810_33_fu_16341_p2[34:14]}};

assign trunc_ln818_54_fu_14386_p4 = {{grp_fu_21752_p2[28:14]}};

assign trunc_ln818_55_fu_16546_p4 = {{add_ln810_34_fu_16532_p2[34:14]}};

assign trunc_ln818_56_fu_14560_p4 = {{grp_fu_21764_p2[33:14]}};

assign trunc_ln818_57_fu_16716_p4 = {{add_ln810_35_fu_16703_p2[34:14]}};

assign trunc_ln818_58_fu_18172_p4 = {{add_ln810_36_fu_18159_p2[34:14]}};

assign trunc_ln818_59_fu_14757_p4 = {{grp_fu_21783_p2[29:14]}};

assign trunc_ln818_5_fu_5319_p4 = {{add_ln810_4_fu_5305_p2[34:14]}};

assign trunc_ln818_60_fu_16953_p4 = {{add_ln810_37_fu_16939_p2[34:14]}};

assign trunc_ln818_61_fu_18384_p4 = {{add_ln810_38_fu_18370_p2[34:14]}};

assign trunc_ln818_62_fu_12656_p4 = {{sub_ln1273_6_fu_12642_p2[34:14]}};

assign trunc_ln818_63_fu_12877_p4 = {{sub_ln1273_7_fu_12863_p2[34:14]}};

assign trunc_ln818_64_fu_13026_p4 = {{sub_ln1273_8_fu_13012_p2[34:14]}};

assign trunc_ln818_6_fu_6009_p4 = {{add_ln810_5_fu_5996_p2[34:14]}};

assign trunc_ln818_7_fu_6705_p4 = {{add_ln810_6_fu_6691_p2[34:14]}};

assign trunc_ln818_8_fu_7417_p4 = {{add_ln810_7_fu_7404_p2[34:14]}};

assign trunc_ln818_9_fu_8201_p4 = {{add_ln810_8_fu_8187_p2[34:14]}};

assign trunc_ln818_s_fu_8824_p4 = {{add_ln810_9_fu_8810_p2[34:14]}};

assign trunc_ln_fu_1984_p4 = {{grp_fu_21385_p2[34:14]}};

assign xk_admm_V_0 = select_ln346_139_fu_12187_p3;

assign xor_ln302_10_fu_2979_p2 = (tmp_56_fu_2959_p3 ^ tmp_55_fu_2945_p3);

assign xor_ln302_11_fu_3049_p2 = (tmp_58_fu_3029_p3 ^ tmp_57_fu_3015_p3);

assign xor_ln302_12_fu_3698_p2 = (tmp_60_fu_3678_p3 ^ tmp_59_fu_3664_p3);

assign xor_ln302_13_fu_3768_p2 = (tmp_62_fu_3748_p3 ^ tmp_61_fu_3734_p3);

assign xor_ln302_14_fu_4555_p2 = (tmp_64_fu_4535_p3 ^ tmp_63_fu_4521_p3);

assign xor_ln302_15_fu_4625_p2 = (tmp_66_fu_4605_p3 ^ tmp_65_fu_4591_p3);

assign xor_ln302_16_fu_5190_p2 = (tmp_68_fu_5170_p3 ^ tmp_67_fu_5156_p3);

assign xor_ln302_17_fu_5260_p2 = (tmp_70_fu_5240_p3 ^ tmp_69_fu_5226_p3);

assign xor_ln302_18_fu_1427_p2 = (tmp_38_fu_1407_p3 ^ tmp_37_fu_1393_p3);

assign xor_ln302_19_fu_1505_p2 = (tmp_40_fu_1485_p3 ^ tmp_39_fu_1471_p3);

assign xor_ln302_20_fu_1657_p2 = (tmp_42_fu_1637_p3 ^ tmp_41_fu_1623_p3);

assign xor_ln302_21_fu_10318_p2 = (tmp_288_fu_10298_p3 ^ tmp_287_fu_10286_p3);

assign xor_ln302_22_fu_9596_p2 = (tmp_290_fu_9576_p3 ^ tmp_289_fu_9564_p3);

assign xor_ln302_23_fu_8695_p2 = (tmp_292_fu_8675_p3 ^ tmp_291_fu_8663_p3);

assign xor_ln302_24_fu_18607_p2 = (tmp_545_fu_18587_p3 ^ tmp_544_fu_18573_p3);

assign xor_ln302_25_fu_18678_p2 = (tmp_547_fu_18658_p3 ^ tmp_546_fu_18644_p3);

assign xor_ln302_26_fu_18783_p2 = (tmp_549_fu_18763_p3 ^ tmp_548_fu_18749_p3);

assign xor_ln302_27_fu_18854_p2 = (tmp_551_fu_18834_p3 ^ tmp_550_fu_18820_p3);

assign xor_ln302_28_fu_18959_p2 = (tmp_553_fu_18939_p3 ^ tmp_552_fu_18925_p3);

assign xor_ln302_29_fu_19030_p2 = (tmp_555_fu_19010_p3 ^ tmp_554_fu_18996_p3);

assign xor_ln302_30_fu_19135_p2 = (tmp_557_fu_19115_p3 ^ tmp_556_fu_19101_p3);

assign xor_ln302_31_fu_19206_p2 = (tmp_559_fu_19186_p3 ^ tmp_558_fu_19172_p3);

assign xor_ln302_32_fu_19311_p2 = (tmp_561_fu_19291_p3 ^ tmp_560_fu_19277_p3);

assign xor_ln302_33_fu_19382_p2 = (tmp_563_fu_19362_p3 ^ tmp_562_fu_19348_p3);

assign xor_ln302_34_fu_19487_p2 = (tmp_565_fu_19467_p3 ^ tmp_564_fu_19453_p3);

assign xor_ln302_35_fu_19558_p2 = (tmp_567_fu_19538_p3 ^ tmp_566_fu_19524_p3);

assign xor_ln302_36_fu_19663_p2 = (tmp_569_fu_19643_p3 ^ tmp_568_fu_19629_p3);

assign xor_ln302_37_fu_19734_p2 = (tmp_571_fu_19714_p3 ^ tmp_570_fu_19700_p3);

assign xor_ln302_38_fu_19839_p2 = (tmp_573_fu_19819_p3 ^ tmp_572_fu_19805_p3);

assign xor_ln302_39_fu_19910_p2 = (tmp_575_fu_19890_p3 ^ tmp_574_fu_19876_p3);

assign xor_ln302_40_fu_20015_p2 = (tmp_577_fu_19995_p3 ^ tmp_576_fu_19981_p3);

assign xor_ln302_41_fu_20086_p2 = (tmp_579_fu_20066_p3 ^ tmp_578_fu_20052_p3);

assign xor_ln302_42_fu_20189_p2 = (tmp_581_fu_20169_p3 ^ tmp_580_fu_20156_p3);

assign xor_ln302_43_fu_20258_p2 = (tmp_583_fu_20238_p3 ^ tmp_582_fu_20225_p3);

assign xor_ln302_44_fu_20327_p2 = (tmp_585_fu_20307_p3 ^ tmp_584_fu_20294_p3);

assign xor_ln302_45_fu_20396_p2 = (tmp_587_fu_20376_p3 ^ tmp_586_fu_20363_p3);

assign xor_ln302_46_fu_20465_p2 = (tmp_589_fu_20445_p3 ^ tmp_588_fu_20432_p3);

assign xor_ln302_47_fu_20534_p2 = (tmp_591_fu_20514_p3 ^ tmp_590_fu_20501_p3);

assign xor_ln302_48_fu_20603_p2 = (tmp_593_fu_20583_p3 ^ tmp_592_fu_20570_p3);

assign xor_ln302_49_fu_20672_p2 = (tmp_595_fu_20652_p3 ^ tmp_594_fu_20639_p3);

assign xor_ln302_4_fu_1575_p2 = (tmp_44_fu_1555_p3 ^ tmp_43_fu_1541_p3);

assign xor_ln302_50_fu_20741_p2 = (tmp_597_fu_20721_p3 ^ tmp_596_fu_20708_p3);

assign xor_ln302_51_fu_20810_p2 = (tmp_599_fu_20790_p3 ^ tmp_598_fu_20777_p3);

assign xor_ln302_52_fu_20879_p2 = (tmp_601_fu_20859_p3 ^ tmp_600_fu_20846_p3);

assign xor_ln302_53_fu_20948_p2 = (tmp_603_fu_20928_p3 ^ tmp_602_fu_20915_p3);

assign xor_ln302_54_fu_21017_p2 = (tmp_605_fu_20997_p3 ^ tmp_604_fu_20984_p3);

assign xor_ln302_55_fu_21086_p2 = (tmp_607_fu_21066_p3 ^ tmp_606_fu_21053_p3);

assign xor_ln302_56_fu_21155_p2 = (tmp_609_fu_21135_p3 ^ tmp_608_fu_21122_p3);

assign xor_ln302_57_fu_21224_p2 = (tmp_611_fu_21204_p3 ^ tmp_610_fu_21191_p3);

assign xor_ln302_58_fu_21293_p2 = (tmp_613_fu_21273_p3 ^ tmp_612_fu_21260_p3);

assign xor_ln302_59_fu_21362_p2 = (tmp_615_fu_21342_p3 ^ tmp_614_fu_21329_p3);

assign xor_ln302_5_fu_1727_p2 = (tmp_46_fu_1707_p3 ^ tmp_45_fu_1693_p3);

assign xor_ln302_6_fu_1885_p2 = (tmp_48_fu_1865_p3 ^ tmp_47_fu_1851_p3);

assign xor_ln302_7_fu_1955_p2 = (tmp_50_fu_1935_p3 ^ tmp_49_fu_1921_p3);

assign xor_ln302_8_fu_2226_p2 = (tmp_52_fu_2206_p3 ^ tmp_51_fu_2192_p3);

assign xor_ln302_9_fu_2296_p2 = (tmp_54_fu_2276_p3 ^ tmp_53_fu_2262_p3);

assign xor_ln302_fu_1357_p2 = (tmp_fu_1323_p3 ^ tmp_36_fu_1337_p3);

assign xor_ln346_10_fu_4343_p2 = (tmp_248_fu_4315_p3 ^ tmp_247_fu_4307_p3);

assign xor_ln346_11_fu_4393_p2 = (tmp_250_fu_4365_p3 ^ tmp_249_fu_4357_p3);

assign xor_ln346_12_fu_4443_p2 = (tmp_252_fu_4415_p3 ^ tmp_251_fu_4407_p3);

assign xor_ln346_13_fu_4485_p2 = (tmp_254_fu_4465_p3 ^ tmp_253_fu_4457_p3);

assign xor_ln346_14_fu_7158_p2 = (tmp_268_fu_7130_p3 ^ tmp_267_fu_7122_p3);

assign xor_ln346_15_fu_7200_p2 = (tmp_270_fu_7180_p3 ^ tmp_269_fu_7172_p3);

assign xor_ln346_16_fu_7908_p2 = (tmp_278_fu_7880_p3 ^ tmp_277_fu_7872_p3);

assign xor_ln346_17_fu_7950_p2 = (tmp_280_fu_7930_p3 ^ tmp_279_fu_7922_p3);

assign xor_ln346_18_fu_14980_p2 = (tmp_354_fu_14952_p3 ^ tmp_353_fu_14944_p3);

assign xor_ln346_19_fu_15030_p2 = (tmp_356_fu_15002_p3 ^ tmp_355_fu_14994_p3);

assign xor_ln346_1_fu_9958_p2 = (tmp_152_fu_9938_p3 ^ tmp_151_fu_9930_p3);

assign xor_ln346_20_fu_15098_p2 = (tmp_364_fu_15070_p3 ^ tmp_363_fu_15062_p3);

assign xor_ln346_21_fu_15148_p2 = (tmp_366_fu_15120_p3 ^ tmp_365_fu_15112_p3);

assign xor_ln346_22_fu_17209_p2 = (tmp_380_fu_17181_p3 ^ tmp_379_fu_17173_p3);

assign xor_ln346_23_fu_17297_p2 = (tmp_394_fu_17269_p3 ^ tmp_393_fu_17261_p3);

assign xor_ln346_24_fu_17780_p2 = (tmp_438_fu_17752_p3 ^ tmp_437_fu_17744_p3);

assign xor_ln346_25_fu_17830_p2 = (tmp_440_fu_17802_p3 ^ tmp_439_fu_17794_p3);

assign xor_ln346_26_fu_17898_p2 = (tmp_448_fu_17870_p3 ^ tmp_447_fu_17862_p3);

assign xor_ln346_27_fu_17948_p2 = (tmp_450_fu_17920_p3 ^ tmp_449_fu_17912_p3);

assign xor_ln346_28_fu_18037_p2 = (tmp_464_fu_18009_p3 ^ tmp_463_fu_18001_p3);

assign xor_ln346_29_fu_18125_p2 = (tmp_478_fu_18097_p3 ^ tmp_477_fu_18089_p3);

assign xor_ln346_2_fu_10213_p2 = (tmp_160_fu_10185_p3 ^ tmp_159_fu_10177_p3);

assign xor_ln346_30_fu_12276_p2 = (tmp_516_fu_12248_p3 ^ tmp_515_fu_12240_p3);

assign xor_ln346_31_fu_12326_p2 = (tmp_518_fu_12298_p3 ^ tmp_517_fu_12290_p3);

assign xor_ln346_32_fu_12376_p2 = (tmp_520_fu_12348_p3 ^ tmp_519_fu_12340_p3);

assign xor_ln346_33_fu_12509_p2 = (tmp_525_fu_12481_p3 ^ tmp_524_fu_12473_p3);

assign xor_ln346_34_fu_12776_p2 = (tmp_533_fu_12748_p3 ^ tmp_532_fu_12740_p3);

assign xor_ln346_35_fu_12826_p2 = (tmp_535_fu_12798_p3 ^ tmp_534_fu_12790_p3);

assign xor_ln346_36_fu_12997_p2 = (tmp_540_fu_12969_p3 ^ tmp_539_fu_12961_p3);

assign xor_ln346_3_fu_10263_p2 = (tmp_162_fu_10235_p3 ^ tmp_161_fu_10227_p3);

assign xor_ln346_4_fu_5557_p2 = (tmp_188_fu_5529_p3 ^ tmp_187_fu_5521_p3);

assign xor_ln346_5_fu_5599_p2 = (tmp_190_fu_5579_p3 ^ tmp_189_fu_5571_p3);

assign xor_ln346_6_fu_8410_p2 = (tmp_216_fu_8390_p3 ^ tmp_215_fu_8382_p3);

assign xor_ln346_7_fu_9048_p2 = (tmp_224_fu_9020_p3 ^ tmp_223_fu_9012_p3);

assign xor_ln346_8_fu_9090_p2 = (tmp_226_fu_9070_p3 ^ tmp_225_fu_9062_p3);

assign xor_ln346_9_fu_9541_p2 = (tmp_234_fu_9513_p3 ^ tmp_233_fu_9505_p3);

assign xor_ln346_fu_9916_p2 = (tmp_150_fu_9888_p3 ^ tmp_149_fu_9880_p3);

assign xor_ln888_100_fu_17611_p2 = (tmp_426_fu_17566_p3 ^ 1'd1);

assign xor_ln888_101_fu_17623_p2 = (tmp_429_fu_17603_p3 ^ or_ln888_50_fu_17617_p2);

assign xor_ln888_102_fu_16044_p2 = (tmp_432_fu_15993_p3 ^ 1'd1);

assign xor_ln888_103_fu_16056_p2 = (tmp_435_fu_16037_p3 ^ or_ln888_51_fu_16050_p2);

assign xor_ln888_104_fu_16218_p2 = (tmp_442_fu_16167_p3 ^ 1'd1);

assign xor_ln888_105_fu_16230_p2 = (tmp_445_fu_16211_p3 ^ or_ln888_52_fu_16224_p2);

assign xor_ln888_106_fu_14260_p2 = (tmp_452_fu_14209_p3 ^ 1'd1);

assign xor_ln888_107_fu_14272_p2 = (tmp_455_fu_14253_p3 ^ or_ln888_53_fu_14266_p2);

assign xor_ln888_108_fu_16411_p2 = (tmp_458_fu_16364_p3 ^ 1'd1);

assign xor_ln888_109_fu_16423_p2 = (tmp_461_fu_16403_p3 ^ or_ln888_54_fu_16417_p2);

assign xor_ln888_10_fu_5374_p2 = (tmp_102_fu_5329_p3 ^ 1'd1);

assign xor_ln888_110_fu_14450_p2 = (tmp_466_fu_14399_p3 ^ 1'd1);

assign xor_ln888_111_fu_14462_p2 = (tmp_469_fu_14443_p3 ^ or_ln888_55_fu_14456_p2);

assign xor_ln888_112_fu_16603_p2 = (tmp_472_fu_16556_p3 ^ 1'd1);

assign xor_ln888_113_fu_16615_p2 = (tmp_475_fu_16595_p3 ^ or_ln888_56_fu_16609_p2);

assign xor_ln888_114_fu_14624_p2 = (tmp_480_fu_14573_p3 ^ 1'd1);

assign xor_ln888_115_fu_14636_p2 = (tmp_483_fu_14617_p3 ^ or_ln888_57_fu_14630_p2);

assign xor_ln888_116_fu_16771_p2 = (tmp_486_fu_16726_p3 ^ 1'd1);

assign xor_ln888_117_fu_16783_p2 = (tmp_489_fu_16763_p3 ^ or_ln888_58_fu_16777_p2);

assign xor_ln888_118_fu_18227_p2 = (tmp_492_fu_18182_p3 ^ 1'd1);

assign xor_ln888_119_fu_18239_p2 = (tmp_495_fu_18219_p3 ^ or_ln888_59_fu_18233_p2);

assign xor_ln888_11_fu_5386_p2 = (tmp_105_fu_5366_p3 ^ or_ln888_5_fu_5380_p2);

assign xor_ln888_120_fu_14821_p2 = (tmp_498_fu_14770_p3 ^ 1'd1);

assign xor_ln888_121_fu_14833_p2 = (tmp_501_fu_14814_p3 ^ or_ln888_60_fu_14827_p2);

assign xor_ln888_122_fu_17008_p2 = (tmp_504_fu_16963_p3 ^ 1'd1);

assign xor_ln888_123_fu_17020_p2 = (tmp_507_fu_17000_p3 ^ or_ln888_61_fu_17014_p2);

assign xor_ln888_124_fu_18439_p2 = (tmp_510_fu_18394_p3 ^ 1'd1);

assign xor_ln888_125_fu_18451_p2 = (tmp_513_fu_18431_p3 ^ or_ln888_62_fu_18445_p2);

assign xor_ln888_12_fu_6064_p2 = (tmp_108_fu_6019_p3 ^ 1'd1);

assign xor_ln888_13_fu_6076_p2 = (tmp_111_fu_6056_p3 ^ or_ln888_6_fu_6070_p2);

assign xor_ln888_14_fu_6760_p2 = (tmp_114_fu_6715_p3 ^ 1'd1);

assign xor_ln888_15_fu_6772_p2 = (tmp_117_fu_6752_p3 ^ or_ln888_7_fu_6766_p2);

assign xor_ln888_16_fu_7472_p2 = (tmp_120_fu_7427_p3 ^ 1'd1);

assign xor_ln888_17_fu_7484_p2 = (tmp_123_fu_7464_p3 ^ or_ln888_8_fu_7478_p2);

assign xor_ln888_18_fu_8265_p2 = (tmp_126_fu_8211_p3 ^ 1'd1);

assign xor_ln888_19_fu_8277_p2 = (tmp_129_fu_8257_p3 ^ or_ln888_9_fu_8271_p2);

assign xor_ln888_1_fu_2056_p2 = (tmp_75_fu_2037_p3 ^ or_ln888_fu_2050_p2);

assign xor_ln888_20_fu_8879_p2 = (tmp_132_fu_8834_p3 ^ 1'd1);

assign xor_ln888_21_fu_8891_p2 = (tmp_135_fu_8871_p3 ^ or_ln888_10_fu_8885_p2);

assign xor_ln888_22_fu_9388_p2 = (tmp_138_fu_9343_p3 ^ 1'd1);

assign xor_ln888_23_fu_9400_p2 = (tmp_141_fu_9380_p3 ^ or_ln888_11_fu_9394_p2);

assign xor_ln888_24_fu_9749_p2 = (tmp_144_fu_9704_p3 ^ 1'd1);

assign xor_ln888_25_fu_9761_p2 = (tmp_147_fu_9741_p3 ^ or_ln888_12_fu_9755_p2);

assign xor_ln888_26_fu_10060_p2 = (tmp_154_fu_10015_p3 ^ 1'd1);

assign xor_ln888_27_fu_10072_p2 = (tmp_157_fu_10052_p3 ^ or_ln888_13_fu_10066_p2);

assign xor_ln888_28_fu_2619_p2 = (tmp_164_fu_2568_p3 ^ 1'd1);

assign xor_ln888_29_fu_2631_p2 = (tmp_167_fu_2612_p3 ^ or_ln888_14_fu_2625_p2);

assign xor_ln888_2_fu_2410_p2 = (tmp_78_fu_2365_p3 ^ 1'd1);

assign xor_ln888_30_fu_3396_p2 = (tmp_170_fu_3349_p3 ^ 1'd1);

assign xor_ln888_31_fu_3408_p2 = (tmp_173_fu_3388_p3 ^ or_ln888_15_fu_3402_p2);

assign xor_ln888_32_fu_4161_p2 = (tmp_176_fu_4116_p3 ^ 1'd1);

assign xor_ln888_33_fu_4173_p2 = (tmp_179_fu_4153_p3 ^ or_ln888_16_fu_4167_p2);

assign xor_ln888_34_fu_5020_p2 = (tmp_182_fu_4975_p3 ^ 1'd1);

assign xor_ln888_35_fu_5032_p2 = (tmp_185_fu_5012_p3 ^ or_ln888_17_fu_5026_p2);

assign xor_ln888_36_fu_5704_p2 = (tmp_192_fu_5665_p3 ^ 1'd1);

assign xor_ln888_37_fu_5716_p2 = (tmp_195_fu_5696_p3 ^ or_ln888_18_fu_5710_p2);

assign xor_ln888_38_fu_6322_p2 = (tmp_198_fu_6277_p3 ^ 1'd1);

assign xor_ln888_39_fu_6334_p2 = (tmp_201_fu_6314_p3 ^ or_ln888_19_fu_6328_p2);

assign xor_ln888_3_fu_2422_p2 = (tmp_81_fu_2402_p3 ^ or_ln888_1_fu_2416_p2);

assign xor_ln888_40_fu_6989_p2 = (tmp_204_fu_6944_p3 ^ 1'd1);

assign xor_ln888_41_fu_7001_p2 = (tmp_207_fu_6981_p3 ^ or_ln888_20_fu_6995_p2);

assign xor_ln888_42_fu_7723_p2 = (tmp_210_fu_7669_p3 ^ 1'd1);

assign xor_ln888_43_fu_7735_p2 = (tmp_213_fu_7715_p3 ^ or_ln888_21_fu_7729_p2);

assign xor_ln888_44_fu_8512_p2 = (tmp_218_fu_8467_p3 ^ 1'd1);

assign xor_ln888_45_fu_8524_p2 = (tmp_221_fu_8504_p3 ^ or_ln888_22_fu_8518_p2);

assign xor_ln888_46_fu_9192_p2 = (tmp_228_fu_9147_p3 ^ 1'd1);

assign xor_ln888_47_fu_9204_p2 = (tmp_231_fu_9184_p3 ^ or_ln888_23_fu_9198_p2);

assign xor_ln888_48_fu_2812_p2 = (tmp_236_fu_2761_p3 ^ 1'd1);

assign xor_ln888_49_fu_2824_p2 = (tmp_239_fu_2805_p3 ^ or_ln888_24_fu_2818_p2);

assign xor_ln888_4_fu_3159_p2 = (tmp_84_fu_3114_p3 ^ 1'd1);

assign xor_ln888_50_fu_3570_p2 = (tmp_242_fu_3523_p3 ^ 1'd1);

assign xor_ln888_51_fu_3582_p2 = (tmp_245_fu_3562_p3 ^ or_ln888_25_fu_3576_p2);

assign xor_ln888_52_fu_5885_p2 = (tmp_256_fu_5838_p3 ^ 1'd1);

assign xor_ln888_53_fu_5897_p2 = (tmp_259_fu_5877_p3 ^ or_ln888_26_fu_5891_p2);

assign xor_ln888_54_fu_6564_p2 = (tmp_262_fu_6519_p3 ^ 1'd1);

assign xor_ln888_55_fu_6576_p2 = (tmp_265_fu_6556_p3 ^ or_ln888_27_fu_6570_p2);

assign xor_ln888_56_fu_7304_p2 = (tmp_272_fu_7257_p3 ^ 1'd1);

assign xor_ln888_57_fu_7316_p2 = (tmp_275_fu_7296_p3 ^ or_ln888_28_fu_7310_p2);

assign xor_ln888_58_fu_8054_p2 = (tmp_282_fu_8007_p3 ^ 1'd1);

assign xor_ln888_59_fu_8066_p2 = (tmp_285_fu_8046_p3 ^ or_ln888_29_fu_8060_p2);

assign xor_ln888_5_fu_3171_p2 = (tmp_87_fu_3151_p3 ^ or_ln888_2_fu_3165_p2);

assign xor_ln888_60_fu_10437_p2 = (tmp_294_fu_10386_p3 ^ 1'd1);

assign xor_ln888_61_fu_10449_p2 = (tmp_297_fu_10430_p3 ^ or_ln888_30_fu_10443_p2);

assign xor_ln888_62_fu_10999_p2 = (tmp_300_fu_10954_p3 ^ 1'd1);

assign xor_ln888_63_fu_11011_p2 = (tmp_303_fu_10991_p3 ^ or_ln888_31_fu_11005_p2);

assign xor_ln888_64_fu_11674_p2 = (tmp_306_fu_11629_p3 ^ 1'd1);

assign xor_ln888_65_fu_11686_p2 = (tmp_309_fu_11666_p3 ^ or_ln888_32_fu_11680_p2);

assign xor_ln888_66_fu_10627_p2 = (tmp_312_fu_10576_p3 ^ 1'd1);

assign xor_ln888_67_fu_10639_p2 = (tmp_315_fu_10620_p3 ^ or_ln888_33_fu_10633_p2);

assign xor_ln888_68_fu_11229_p2 = (tmp_318_fu_11184_p3 ^ 1'd1);

assign xor_ln888_69_fu_11241_p2 = (tmp_321_fu_11221_p3 ^ or_ln888_34_fu_11235_p2);

assign xor_ln888_6_fu_3912_p2 = (tmp_90_fu_3867_p3 ^ 1'd1);

assign xor_ln888_70_fu_11870_p2 = (tmp_324_fu_11825_p3 ^ 1'd1);

assign xor_ln888_71_fu_11882_p2 = (tmp_327_fu_11862_p3 ^ or_ln888_35_fu_11876_p2);

assign xor_ln888_72_fu_10801_p2 = (tmp_330_fu_10750_p3 ^ 1'd1);

assign xor_ln888_73_fu_10813_p2 = (tmp_333_fu_10794_p3 ^ or_ln888_36_fu_10807_p2);

assign xor_ln888_74_fu_11478_p2 = (tmp_336_fu_11433_p3 ^ 1'd1);

assign xor_ln888_75_fu_11490_p2 = (tmp_339_fu_11470_p3 ^ or_ln888_37_fu_11484_p2);

assign xor_ln888_76_fu_12076_p2 = (tmp_342_fu_12031_p3 ^ 1'd1);

assign xor_ln888_77_fu_12088_p2 = (tmp_345_fu_12068_p3 ^ or_ln888_38_fu_12082_p2);

assign xor_ln888_78_fu_13178_p2 = (tmp_348_fu_13127_p3 ^ 1'd1);

assign xor_ln888_79_fu_13190_p2 = (tmp_351_fu_13171_p3 ^ or_ln888_39_fu_13184_p2);

assign xor_ln888_7_fu_3924_p2 = (tmp_93_fu_3904_p3 ^ or_ln888_3_fu_3918_p2);

assign xor_ln888_80_fu_13352_p2 = (tmp_358_fu_13301_p3 ^ 1'd1);

assign xor_ln888_81_fu_13364_p2 = (tmp_361_fu_13345_p3 ^ or_ln888_40_fu_13358_p2);

assign xor_ln888_82_fu_13522_p2 = (tmp_368_fu_13471_p3 ^ 1'd1);

assign xor_ln888_83_fu_13534_p2 = (tmp_371_fu_13515_p3 ^ or_ln888_41_fu_13528_p2);

assign xor_ln888_84_fu_15253_p2 = (tmp_374_fu_15206_p3 ^ 1'd1);

assign xor_ln888_85_fu_15265_p2 = (tmp_377_fu_15245_p3 ^ or_ln888_42_fu_15259_p2);

assign xor_ln888_86_fu_13712_p2 = (tmp_382_fu_13661_p3 ^ 1'd1);

assign xor_ln888_87_fu_13724_p2 = (tmp_385_fu_13705_p3 ^ or_ln888_43_fu_13718_p2);

assign xor_ln888_88_fu_15445_p2 = (tmp_388_fu_15398_p3 ^ 1'd1);

assign xor_ln888_89_fu_15457_p2 = (tmp_391_fu_15437_p3 ^ or_ln888_44_fu_15451_p2);

assign xor_ln888_8_fu_4753_p2 = (tmp_96_fu_4708_p3 ^ 1'd1);

assign xor_ln888_90_fu_13886_p2 = (tmp_396_fu_13835_p3 ^ 1'd1);

assign xor_ln888_91_fu_13898_p2 = (tmp_399_fu_13879_p3 ^ or_ln888_45_fu_13892_p2);

assign xor_ln888_92_fu_15613_p2 = (tmp_402_fu_15568_p3 ^ 1'd1);

assign xor_ln888_93_fu_15625_p2 = (tmp_405_fu_15605_p3 ^ or_ln888_46_fu_15619_p2);

assign xor_ln888_94_fu_17399_p2 = (tmp_408_fu_17354_p3 ^ 1'd1);

assign xor_ln888_95_fu_17411_p2 = (tmp_411_fu_17391_p3 ^ or_ln888_47_fu_17405_p2);

assign xor_ln888_96_fu_14083_p2 = (tmp_414_fu_14032_p3 ^ 1'd1);

assign xor_ln888_97_fu_14095_p2 = (tmp_417_fu_14076_p3 ^ or_ln888_48_fu_14089_p2);

assign xor_ln888_98_fu_15850_p2 = (tmp_420_fu_15805_p3 ^ 1'd1);

assign xor_ln888_99_fu_15862_p2 = (tmp_423_fu_15842_p3 ^ or_ln888_49_fu_15856_p2);

assign xor_ln888_9_fu_4765_p2 = (tmp_99_fu_4745_p3 ^ or_ln888_4_fu_4759_p2);

assign xor_ln888_fu_2044_p2 = (tmp_72_fu_1993_p3 ^ 1'd1);

assign xor_ln890_10_fu_8905_p2 = (tmp_136_fu_8897_p3 ^ 1'd1);

assign xor_ln890_11_fu_9414_p2 = (tmp_142_fu_9406_p3 ^ 1'd1);

assign xor_ln890_12_fu_9775_p2 = (tmp_148_fu_9767_p3 ^ 1'd1);

assign xor_ln890_13_fu_10086_p2 = (tmp_158_fu_10078_p3 ^ 1'd1);

assign xor_ln890_14_fu_2644_p2 = (tmp_168_fu_2637_p3 ^ 1'd1);

assign xor_ln890_15_fu_3422_p2 = (tmp_174_fu_3414_p3 ^ 1'd1);

assign xor_ln890_16_fu_4187_p2 = (tmp_180_fu_4179_p3 ^ 1'd1);

assign xor_ln890_17_fu_5046_p2 = (tmp_186_fu_5038_p3 ^ 1'd1);

assign xor_ln890_18_fu_5730_p2 = (tmp_196_fu_5722_p3 ^ 1'd1);

assign xor_ln890_19_fu_6348_p2 = (tmp_202_fu_6340_p3 ^ 1'd1);

assign xor_ln890_1_fu_2436_p2 = (tmp_82_fu_2428_p3 ^ 1'd1);

assign xor_ln890_20_fu_7015_p2 = (tmp_208_fu_7007_p3 ^ 1'd1);

assign xor_ln890_21_fu_7749_p2 = (tmp_214_fu_7741_p3 ^ 1'd1);

assign xor_ln890_22_fu_8538_p2 = (tmp_222_fu_8530_p3 ^ 1'd1);

assign xor_ln890_23_fu_9218_p2 = (tmp_232_fu_9210_p3 ^ 1'd1);

assign xor_ln890_24_fu_2837_p2 = (tmp_240_fu_2830_p3 ^ 1'd1);

assign xor_ln890_25_fu_3596_p2 = (tmp_246_fu_3588_p3 ^ 1'd1);

assign xor_ln890_26_fu_5911_p2 = (tmp_260_fu_5903_p3 ^ 1'd1);

assign xor_ln890_27_fu_6590_p2 = (tmp_266_fu_6582_p3 ^ 1'd1);

assign xor_ln890_28_fu_7330_p2 = (tmp_276_fu_7322_p3 ^ 1'd1);

assign xor_ln890_29_fu_8080_p2 = (tmp_286_fu_8072_p3 ^ 1'd1);

assign xor_ln890_2_fu_3185_p2 = (tmp_88_fu_3177_p3 ^ 1'd1);

assign xor_ln890_30_fu_10462_p2 = (tmp_298_fu_10455_p3 ^ 1'd1);

assign xor_ln890_31_fu_11025_p2 = (tmp_304_fu_11017_p3 ^ 1'd1);

assign xor_ln890_32_fu_11700_p2 = (tmp_310_fu_11692_p3 ^ 1'd1);

assign xor_ln890_33_fu_10652_p2 = (tmp_316_fu_10645_p3 ^ 1'd1);

assign xor_ln890_34_fu_11255_p2 = (tmp_322_fu_11247_p3 ^ 1'd1);

assign xor_ln890_35_fu_11896_p2 = (tmp_328_fu_11888_p3 ^ 1'd1);

assign xor_ln890_36_fu_10826_p2 = (tmp_334_fu_10819_p3 ^ 1'd1);

assign xor_ln890_37_fu_11504_p2 = (tmp_340_fu_11496_p3 ^ 1'd1);

assign xor_ln890_38_fu_12102_p2 = (tmp_346_fu_12094_p3 ^ 1'd1);

assign xor_ln890_39_fu_13203_p2 = (tmp_352_fu_13196_p3 ^ 1'd1);

assign xor_ln890_3_fu_3938_p2 = (tmp_94_fu_3930_p3 ^ 1'd1);

assign xor_ln890_40_fu_13377_p2 = (tmp_362_fu_13370_p3 ^ 1'd1);

assign xor_ln890_41_fu_13547_p2 = (tmp_372_fu_13540_p3 ^ 1'd1);

assign xor_ln890_42_fu_15279_p2 = (tmp_378_fu_15271_p3 ^ 1'd1);

assign xor_ln890_43_fu_13737_p2 = (tmp_386_fu_13730_p3 ^ 1'd1);

assign xor_ln890_44_fu_15471_p2 = (tmp_392_fu_15463_p3 ^ 1'd1);

assign xor_ln890_45_fu_13911_p2 = (tmp_400_fu_13904_p3 ^ 1'd1);

assign xor_ln890_46_fu_15639_p2 = (tmp_406_fu_15631_p3 ^ 1'd1);

assign xor_ln890_47_fu_17425_p2 = (tmp_412_fu_17417_p3 ^ 1'd1);

assign xor_ln890_48_fu_14108_p2 = (tmp_418_fu_14101_p3 ^ 1'd1);

assign xor_ln890_49_fu_15876_p2 = (tmp_424_fu_15868_p3 ^ 1'd1);

assign xor_ln890_4_fu_4779_p2 = (tmp_100_fu_4771_p3 ^ 1'd1);

assign xor_ln890_50_fu_17637_p2 = (tmp_430_fu_17629_p3 ^ 1'd1);

assign xor_ln890_51_fu_16069_p2 = (tmp_436_fu_16062_p3 ^ 1'd1);

assign xor_ln890_52_fu_16243_p2 = (tmp_446_fu_16236_p3 ^ 1'd1);

assign xor_ln890_53_fu_14285_p2 = (tmp_456_fu_14278_p3 ^ 1'd1);

assign xor_ln890_54_fu_16437_p2 = (tmp_462_fu_16429_p3 ^ 1'd1);

assign xor_ln890_55_fu_14475_p2 = (tmp_470_fu_14468_p3 ^ 1'd1);

assign xor_ln890_56_fu_16629_p2 = (tmp_476_fu_16621_p3 ^ 1'd1);

assign xor_ln890_57_fu_14649_p2 = (tmp_484_fu_14642_p3 ^ 1'd1);

assign xor_ln890_58_fu_16797_p2 = (tmp_490_fu_16789_p3 ^ 1'd1);

assign xor_ln890_59_fu_18253_p2 = (tmp_496_fu_18245_p3 ^ 1'd1);

assign xor_ln890_5_fu_5400_p2 = (tmp_106_fu_5392_p3 ^ 1'd1);

assign xor_ln890_60_fu_14846_p2 = (tmp_502_fu_14839_p3 ^ 1'd1);

assign xor_ln890_61_fu_17034_p2 = (tmp_508_fu_17026_p3 ^ 1'd1);

assign xor_ln890_62_fu_18465_p2 = (tmp_514_fu_18457_p3 ^ 1'd1);

assign xor_ln890_6_fu_6090_p2 = (tmp_112_fu_6082_p3 ^ 1'd1);

assign xor_ln890_7_fu_6786_p2 = (tmp_118_fu_6778_p3 ^ 1'd1);

assign xor_ln890_8_fu_7498_p2 = (tmp_124_fu_7490_p3 ^ 1'd1);

assign xor_ln890_9_fu_8291_p2 = (tmp_130_fu_8283_p3 ^ 1'd1);

assign xor_ln890_fu_2069_p2 = (tmp_76_fu_2062_p3 ^ 1'd1);

assign xor_ln895_100_fu_7360_p2 = (tmp_271_fu_7239_p3 ^ 1'd1);

assign xor_ln895_101_fu_7888_p2 = (tmp_277_fu_7872_p3 ^ 1'd1);

assign xor_ln895_102_fu_7938_p2 = (tmp_279_fu_7922_p3 ^ 1'd1);

assign xor_ln895_103_fu_8098_p2 = (xor_ln888_59_fu_8066_p2 ^ 1'd1);

assign xor_ln895_104_fu_8110_p2 = (tmp_281_fu_7989_p3 ^ 1'd1);

assign xor_ln895_105_fu_10306_p2 = (tmp_287_fu_10286_p3 ^ 1'd1);

assign xor_ln895_106_fu_9584_p2 = (tmp_289_fu_9564_p3 ^ 1'd1);

assign xor_ln895_107_fu_8683_p2 = (tmp_291_fu_8663_p3 ^ 1'd1);

assign xor_ln895_108_fu_10486_p2 = (xor_ln888_61_fu_10449_p2 ^ 1'd1);

assign xor_ln895_109_fu_10498_p2 = (tmp_293_fu_10366_p3 ^ 1'd1);

assign xor_ln895_10_fu_2967_p2 = (tmp_55_fu_2945_p3 ^ 1'd1);

assign xor_ln895_110_fu_11049_p2 = (xor_ln888_63_fu_11011_p2 ^ 1'd1);

assign xor_ln895_111_fu_11061_p2 = (tmp_299_fu_10936_p3 ^ 1'd1);

assign xor_ln895_112_fu_11724_p2 = (xor_ln888_65_fu_11686_p2 ^ 1'd1);

assign xor_ln895_113_fu_11736_p2 = (tmp_305_fu_11611_p3 ^ 1'd1);

assign xor_ln895_114_fu_10676_p2 = (xor_ln888_67_fu_10639_p2 ^ 1'd1);

assign xor_ln895_115_fu_10688_p2 = (tmp_311_fu_10556_p3 ^ 1'd1);

assign xor_ln895_116_fu_11279_p2 = (xor_ln888_69_fu_11241_p2 ^ 1'd1);

assign xor_ln895_117_fu_11291_p2 = (tmp_317_fu_11166_p3 ^ 1'd1);

assign xor_ln895_118_fu_11920_p2 = (xor_ln888_71_fu_11882_p2 ^ 1'd1);

assign xor_ln895_119_fu_11932_p2 = (tmp_323_fu_11807_p3 ^ 1'd1);

assign xor_ln895_11_fu_3037_p2 = (tmp_57_fu_3015_p3 ^ 1'd1);

assign xor_ln895_120_fu_10850_p2 = (xor_ln888_73_fu_10813_p2 ^ 1'd1);

assign xor_ln895_121_fu_10862_p2 = (tmp_329_fu_10730_p3 ^ 1'd1);

assign xor_ln895_122_fu_11528_p2 = (xor_ln888_75_fu_11490_p2 ^ 1'd1);

assign xor_ln895_123_fu_11540_p2 = (tmp_335_fu_11415_p3 ^ 1'd1);

assign xor_ln895_124_fu_12126_p2 = (xor_ln888_77_fu_12088_p2 ^ 1'd1);

assign xor_ln895_125_fu_12138_p2 = (tmp_341_fu_12013_p3 ^ 1'd1);

assign xor_ln895_126_fu_13227_p2 = (xor_ln888_79_fu_13190_p2 ^ 1'd1);

assign xor_ln895_127_fu_13239_p2 = (tmp_347_fu_13111_p3 ^ 1'd1);

assign xor_ln895_128_fu_14960_p2 = (tmp_353_fu_14944_p3 ^ 1'd1);

assign xor_ln895_129_fu_15010_p2 = (tmp_355_fu_14994_p3 ^ 1'd1);

assign xor_ln895_12_fu_3686_p2 = (tmp_59_fu_3664_p3 ^ 1'd1);

assign xor_ln895_130_fu_13401_p2 = (xor_ln888_81_fu_13364_p2 ^ 1'd1);

assign xor_ln895_131_fu_13413_p2 = (tmp_357_fu_13281_p3 ^ 1'd1);

assign xor_ln895_132_fu_15078_p2 = (tmp_363_fu_15062_p3 ^ 1'd1);

assign xor_ln895_133_fu_15128_p2 = (tmp_365_fu_15112_p3 ^ 1'd1);

assign xor_ln895_134_fu_13571_p2 = (xor_ln888_83_fu_13534_p2 ^ 1'd1);

assign xor_ln895_135_fu_13583_p2 = (tmp_367_fu_13455_p3 ^ 1'd1);

assign xor_ln895_136_fu_15297_p2 = (xor_ln888_85_fu_15265_p2 ^ 1'd1);

assign xor_ln895_137_fu_15309_p2 = (tmp_373_fu_15188_p3 ^ 1'd1);

assign xor_ln895_138_fu_17189_p2 = (tmp_379_fu_17173_p3 ^ 1'd1);

assign xor_ln895_139_fu_13761_p2 = (xor_ln888_87_fu_13724_p2 ^ 1'd1);

assign xor_ln895_13_fu_3756_p2 = (tmp_61_fu_3734_p3 ^ 1'd1);

assign xor_ln895_140_fu_13773_p2 = (tmp_381_fu_13641_p3 ^ 1'd1);

assign xor_ln895_141_fu_15489_p2 = (xor_ln888_89_fu_15457_p2 ^ 1'd1);

assign xor_ln895_142_fu_15501_p2 = (tmp_387_fu_15380_p3 ^ 1'd1);

assign xor_ln895_143_fu_17277_p2 = (tmp_393_fu_17261_p3 ^ 1'd1);

assign xor_ln895_144_fu_13935_p2 = (xor_ln888_91_fu_13898_p2 ^ 1'd1);

assign xor_ln895_145_fu_13947_p2 = (tmp_395_fu_13815_p3 ^ 1'd1);

assign xor_ln895_146_fu_15663_p2 = (xor_ln888_93_fu_15625_p2 ^ 1'd1);

assign xor_ln895_147_fu_15675_p2 = (tmp_401_fu_15550_p3 ^ 1'd1);

assign xor_ln895_148_fu_17449_p2 = (xor_ln888_95_fu_17411_p2 ^ 1'd1);

assign xor_ln895_149_fu_17461_p2 = (tmp_407_fu_17336_p3 ^ 1'd1);

assign xor_ln895_14_fu_4543_p2 = (tmp_63_fu_4521_p3 ^ 1'd1);

assign xor_ln895_150_fu_14132_p2 = (xor_ln888_97_fu_14095_p2 ^ 1'd1);

assign xor_ln895_151_fu_14144_p2 = (tmp_413_fu_14012_p3 ^ 1'd1);

assign xor_ln895_152_fu_15900_p2 = (xor_ln888_99_fu_15862_p2 ^ 1'd1);

assign xor_ln895_153_fu_15912_p2 = (tmp_419_fu_15787_p3 ^ 1'd1);

assign xor_ln895_154_fu_17661_p2 = (xor_ln888_101_fu_17623_p2 ^ 1'd1);

assign xor_ln895_155_fu_17673_p2 = (tmp_425_fu_17548_p3 ^ 1'd1);

assign xor_ln895_156_fu_16093_p2 = (xor_ln888_103_fu_16056_p2 ^ 1'd1);

assign xor_ln895_157_fu_16105_p2 = (tmp_431_fu_15977_p3 ^ 1'd1);

assign xor_ln895_158_fu_17760_p2 = (tmp_437_fu_17744_p3 ^ 1'd1);

assign xor_ln895_159_fu_17810_p2 = (tmp_439_fu_17794_p3 ^ 1'd1);

assign xor_ln895_15_fu_4613_p2 = (tmp_65_fu_4591_p3 ^ 1'd1);

assign xor_ln895_160_fu_16267_p2 = (xor_ln888_105_fu_16230_p2 ^ 1'd1);

assign xor_ln895_161_fu_16279_p2 = (tmp_441_fu_16147_p3 ^ 1'd1);

assign xor_ln895_162_fu_17878_p2 = (tmp_447_fu_17862_p3 ^ 1'd1);

assign xor_ln895_163_fu_17928_p2 = (tmp_449_fu_17912_p3 ^ 1'd1);

assign xor_ln895_164_fu_14309_p2 = (xor_ln888_107_fu_14272_p2 ^ 1'd1);

assign xor_ln895_165_fu_14321_p2 = (tmp_451_fu_14193_p3 ^ 1'd1);

assign xor_ln895_166_fu_16455_p2 = (xor_ln888_109_fu_16423_p2 ^ 1'd1);

assign xor_ln895_167_fu_16467_p2 = (tmp_457_fu_16346_p3 ^ 1'd1);

assign xor_ln895_168_fu_18017_p2 = (tmp_463_fu_18001_p3 ^ 1'd1);

assign xor_ln895_169_fu_14499_p2 = (xor_ln888_111_fu_14462_p2 ^ 1'd1);

assign xor_ln895_16_fu_5178_p2 = (tmp_67_fu_5156_p3 ^ 1'd1);

assign xor_ln895_170_fu_14511_p2 = (tmp_465_fu_14379_p3 ^ 1'd1);

assign xor_ln895_171_fu_16647_p2 = (xor_ln888_113_fu_16615_p2 ^ 1'd1);

assign xor_ln895_172_fu_16659_p2 = (tmp_471_fu_16538_p3 ^ 1'd1);

assign xor_ln895_173_fu_18105_p2 = (tmp_477_fu_18089_p3 ^ 1'd1);

assign xor_ln895_174_fu_14673_p2 = (xor_ln888_115_fu_14636_p2 ^ 1'd1);

assign xor_ln895_175_fu_14685_p2 = (tmp_479_fu_14553_p3 ^ 1'd1);

assign xor_ln895_176_fu_16821_p2 = (xor_ln888_117_fu_16783_p2 ^ 1'd1);

assign xor_ln895_177_fu_16833_p2 = (tmp_485_fu_16708_p3 ^ 1'd1);

assign xor_ln895_178_fu_18277_p2 = (xor_ln888_119_fu_18239_p2 ^ 1'd1);

assign xor_ln895_179_fu_18289_p2 = (tmp_491_fu_18164_p3 ^ 1'd1);

assign xor_ln895_17_fu_5248_p2 = (tmp_69_fu_5226_p3 ^ 1'd1);

assign xor_ln895_180_fu_14870_p2 = (xor_ln888_121_fu_14833_p2 ^ 1'd1);

assign xor_ln895_181_fu_14882_p2 = (tmp_497_fu_14750_p3 ^ 1'd1);

assign xor_ln895_182_fu_17058_p2 = (xor_ln888_123_fu_17020_p2 ^ 1'd1);

assign xor_ln895_183_fu_17070_p2 = (tmp_503_fu_16945_p3 ^ 1'd1);

assign xor_ln895_184_fu_18489_p2 = (xor_ln888_125_fu_18451_p2 ^ 1'd1);

assign xor_ln895_185_fu_18501_p2 = (tmp_509_fu_18376_p3 ^ 1'd1);

assign xor_ln895_186_fu_12256_p2 = (tmp_515_fu_12240_p3 ^ 1'd1);

assign xor_ln895_187_fu_12306_p2 = (tmp_517_fu_12290_p3 ^ 1'd1);

assign xor_ln895_188_fu_12356_p2 = (tmp_519_fu_12340_p3 ^ 1'd1);

assign xor_ln895_189_fu_12421_p2 = (tmp_521_fu_12391_p3 ^ 1'd1);

assign xor_ln895_18_fu_1415_p2 = (tmp_37_fu_1393_p3 ^ 1'd1);

assign xor_ln895_190_fu_12489_p2 = (tmp_524_fu_12473_p3 ^ 1'd1);

assign xor_ln895_191_fu_12578_p2 = (tmp_526_fu_12548_p3 ^ 1'd1);

assign xor_ln895_192_fu_12688_p2 = (tmp_529_fu_12648_p3 ^ 1'd1);

assign xor_ln895_193_fu_12756_p2 = (tmp_532_fu_12740_p3 ^ 1'd1);

assign xor_ln895_194_fu_12806_p2 = (tmp_534_fu_12790_p3 ^ 1'd1);

assign xor_ln895_195_fu_12909_p2 = (tmp_536_fu_12869_p3 ^ 1'd1);

assign xor_ln895_196_fu_12977_p2 = (tmp_539_fu_12961_p3 ^ 1'd1);

assign xor_ln895_197_fu_13058_p2 = (tmp_541_fu_13018_p3 ^ 1'd1);

assign xor_ln895_198_fu_18595_p2 = (tmp_544_fu_18573_p3 ^ 1'd1);

assign xor_ln895_199_fu_18666_p2 = (tmp_546_fu_18644_p3 ^ 1'd1);

assign xor_ln895_19_fu_1493_p2 = (tmp_39_fu_1471_p3 ^ 1'd1);

assign xor_ln895_200_fu_18771_p2 = (tmp_548_fu_18749_p3 ^ 1'd1);

assign xor_ln895_201_fu_18842_p2 = (tmp_550_fu_18820_p3 ^ 1'd1);

assign xor_ln895_202_fu_18947_p2 = (tmp_552_fu_18925_p3 ^ 1'd1);

assign xor_ln895_203_fu_19018_p2 = (tmp_554_fu_18996_p3 ^ 1'd1);

assign xor_ln895_204_fu_19123_p2 = (tmp_556_fu_19101_p3 ^ 1'd1);

assign xor_ln895_205_fu_19194_p2 = (tmp_558_fu_19172_p3 ^ 1'd1);

assign xor_ln895_206_fu_19299_p2 = (tmp_560_fu_19277_p3 ^ 1'd1);

assign xor_ln895_207_fu_19370_p2 = (tmp_562_fu_19348_p3 ^ 1'd1);

assign xor_ln895_208_fu_19475_p2 = (tmp_564_fu_19453_p3 ^ 1'd1);

assign xor_ln895_209_fu_19546_p2 = (tmp_566_fu_19524_p3 ^ 1'd1);

assign xor_ln895_20_fu_1645_p2 = (tmp_41_fu_1623_p3 ^ 1'd1);

assign xor_ln895_210_fu_19651_p2 = (tmp_568_fu_19629_p3 ^ 1'd1);

assign xor_ln895_211_fu_19722_p2 = (tmp_570_fu_19700_p3 ^ 1'd1);

assign xor_ln895_212_fu_19827_p2 = (tmp_572_fu_19805_p3 ^ 1'd1);

assign xor_ln895_213_fu_19898_p2 = (tmp_574_fu_19876_p3 ^ 1'd1);

assign xor_ln895_214_fu_20003_p2 = (tmp_576_fu_19981_p3 ^ 1'd1);

assign xor_ln895_215_fu_20074_p2 = (tmp_578_fu_20052_p3 ^ 1'd1);

assign xor_ln895_216_fu_20177_p2 = (tmp_580_fu_20156_p3 ^ 1'd1);

assign xor_ln895_217_fu_20246_p2 = (tmp_582_fu_20225_p3 ^ 1'd1);

assign xor_ln895_218_fu_20315_p2 = (tmp_584_fu_20294_p3 ^ 1'd1);

assign xor_ln895_219_fu_20384_p2 = (tmp_586_fu_20363_p3 ^ 1'd1);

assign xor_ln895_21_fu_1563_p2 = (tmp_43_fu_1541_p3 ^ 1'd1);

assign xor_ln895_220_fu_20453_p2 = (tmp_588_fu_20432_p3 ^ 1'd1);

assign xor_ln895_221_fu_20522_p2 = (tmp_590_fu_20501_p3 ^ 1'd1);

assign xor_ln895_222_fu_20591_p2 = (tmp_592_fu_20570_p3 ^ 1'd1);

assign xor_ln895_223_fu_20660_p2 = (tmp_594_fu_20639_p3 ^ 1'd1);

assign xor_ln895_224_fu_20729_p2 = (tmp_596_fu_20708_p3 ^ 1'd1);

assign xor_ln895_225_fu_20798_p2 = (tmp_598_fu_20777_p3 ^ 1'd1);

assign xor_ln895_226_fu_20867_p2 = (tmp_600_fu_20846_p3 ^ 1'd1);

assign xor_ln895_227_fu_20936_p2 = (tmp_602_fu_20915_p3 ^ 1'd1);

assign xor_ln895_228_fu_21005_p2 = (tmp_604_fu_20984_p3 ^ 1'd1);

assign xor_ln895_229_fu_21074_p2 = (tmp_606_fu_21053_p3 ^ 1'd1);

assign xor_ln895_22_fu_1715_p2 = (tmp_45_fu_1693_p3 ^ 1'd1);

assign xor_ln895_230_fu_21143_p2 = (tmp_608_fu_21122_p3 ^ 1'd1);

assign xor_ln895_231_fu_21212_p2 = (tmp_610_fu_21191_p3 ^ 1'd1);

assign xor_ln895_232_fu_21281_p2 = (tmp_612_fu_21260_p3 ^ 1'd1);

assign xor_ln895_233_fu_21350_p2 = (tmp_614_fu_21329_p3 ^ 1'd1);

assign xor_ln895_23_fu_1873_p2 = (tmp_47_fu_1851_p3 ^ 1'd1);

assign xor_ln895_24_fu_1943_p2 = (tmp_49_fu_1921_p3 ^ 1'd1);

assign xor_ln895_25_fu_2214_p2 = (tmp_51_fu_2192_p3 ^ 1'd1);

assign xor_ln895_26_fu_2284_p2 = (tmp_53_fu_2262_p3 ^ 1'd1);

assign xor_ln895_27_fu_2093_p2 = (xor_ln888_1_fu_2056_p2 ^ 1'd1);

assign xor_ln895_28_fu_2105_p2 = (tmp_71_fu_1977_p3 ^ 1'd1);

assign xor_ln895_29_fu_2460_p2 = (xor_ln888_3_fu_2422_p2 ^ 1'd1);

assign xor_ln895_30_fu_2472_p2 = (tmp_77_fu_2347_p3 ^ 1'd1);

assign xor_ln895_31_fu_3209_p2 = (xor_ln888_5_fu_3171_p2 ^ 1'd1);

assign xor_ln895_32_fu_3221_p2 = (tmp_83_fu_3096_p3 ^ 1'd1);

assign xor_ln895_33_fu_3962_p2 = (xor_ln888_7_fu_3924_p2 ^ 1'd1);

assign xor_ln895_34_fu_3974_p2 = (tmp_89_fu_3849_p3 ^ 1'd1);

assign xor_ln895_35_fu_4803_p2 = (xor_ln888_9_fu_4765_p2 ^ 1'd1);

assign xor_ln895_36_fu_4815_p2 = (tmp_95_fu_4690_p3 ^ 1'd1);

assign xor_ln895_37_fu_5424_p2 = (xor_ln888_11_fu_5386_p2 ^ 1'd1);

assign xor_ln895_38_fu_5436_p2 = (tmp_101_fu_5311_p3 ^ 1'd1);

assign xor_ln895_39_fu_6114_p2 = (xor_ln888_13_fu_6076_p2 ^ 1'd1);

assign xor_ln895_40_fu_6126_p2 = (tmp_107_fu_6001_p3 ^ 1'd1);

assign xor_ln895_41_fu_6810_p2 = (xor_ln888_15_fu_6772_p2 ^ 1'd1);

assign xor_ln895_42_fu_6822_p2 = (tmp_113_fu_6697_p3 ^ 1'd1);

assign xor_ln895_43_fu_7522_p2 = (xor_ln888_17_fu_7484_p2 ^ 1'd1);

assign xor_ln895_44_fu_7534_p2 = (tmp_119_fu_7409_p3 ^ 1'd1);

assign xor_ln895_45_fu_8315_p2 = (xor_ln888_19_fu_8277_p2 ^ 1'd1);

assign xor_ln895_46_fu_8327_p2 = (tmp_125_fu_8193_p3 ^ 1'd1);

assign xor_ln895_47_fu_8929_p2 = (xor_ln888_21_fu_8891_p2 ^ 1'd1);

assign xor_ln895_48_fu_8941_p2 = (tmp_131_fu_8816_p3 ^ 1'd1);

assign xor_ln895_49_fu_9438_p2 = (xor_ln888_23_fu_9400_p2 ^ 1'd1);

assign xor_ln895_50_fu_9450_p2 = (tmp_137_fu_9325_p3 ^ 1'd1);

assign xor_ln895_51_fu_9799_p2 = (xor_ln888_25_fu_9761_p2 ^ 1'd1);

assign xor_ln895_52_fu_9811_p2 = (tmp_143_fu_9686_p3 ^ 1'd1);

assign xor_ln895_53_fu_9896_p2 = (tmp_149_fu_9880_p3 ^ 1'd1);

assign xor_ln895_54_fu_9946_p2 = (tmp_151_fu_9930_p3 ^ 1'd1);

assign xor_ln895_55_fu_10110_p2 = (xor_ln888_27_fu_10072_p2 ^ 1'd1);

assign xor_ln895_56_fu_10122_p2 = (tmp_153_fu_9997_p3 ^ 1'd1);

assign xor_ln895_57_fu_10193_p2 = (tmp_159_fu_10177_p3 ^ 1'd1);

assign xor_ln895_58_fu_10243_p2 = (tmp_161_fu_10227_p3 ^ 1'd1);

assign xor_ln895_59_fu_2668_p2 = (xor_ln888_29_fu_2631_p2 ^ 1'd1);

assign xor_ln895_60_fu_2680_p2 = (tmp_163_fu_2552_p3 ^ 1'd1);

assign xor_ln895_61_fu_3440_p2 = (xor_ln888_31_fu_3408_p2 ^ 1'd1);

assign xor_ln895_62_fu_3452_p2 = (tmp_169_fu_3331_p3 ^ 1'd1);

assign xor_ln895_63_fu_4211_p2 = (xor_ln888_33_fu_4173_p2 ^ 1'd1);

assign xor_ln895_64_fu_4223_p2 = (tmp_175_fu_4098_p3 ^ 1'd1);

assign xor_ln895_65_fu_5070_p2 = (xor_ln888_35_fu_5032_p2 ^ 1'd1);

assign xor_ln895_66_fu_5082_p2 = (tmp_181_fu_4957_p3 ^ 1'd1);

assign xor_ln895_67_fu_5537_p2 = (tmp_187_fu_5521_p3 ^ 1'd1);

assign xor_ln895_68_fu_5587_p2 = (tmp_189_fu_5571_p3 ^ 1'd1);

assign xor_ln895_69_fu_5748_p2 = (xor_ln888_37_fu_5716_p2 ^ 1'd1);

assign xor_ln895_70_fu_5760_p2 = (tmp_191_fu_5647_p3 ^ 1'd1);

assign xor_ln895_71_fu_6372_p2 = (xor_ln888_39_fu_6334_p2 ^ 1'd1);

assign xor_ln895_72_fu_6384_p2 = (tmp_197_fu_6259_p3 ^ 1'd1);

assign xor_ln895_73_fu_7039_p2 = (xor_ln888_41_fu_7001_p2 ^ 1'd1);

assign xor_ln895_74_fu_7051_p2 = (tmp_203_fu_6926_p3 ^ 1'd1);

assign xor_ln895_75_fu_7773_p2 = (xor_ln888_43_fu_7735_p2 ^ 1'd1);

assign xor_ln895_76_fu_7785_p2 = (tmp_209_fu_7651_p3 ^ 1'd1);

assign xor_ln895_77_fu_8398_p2 = (tmp_215_fu_8382_p3 ^ 1'd1);

assign xor_ln895_78_fu_8562_p2 = (xor_ln888_45_fu_8524_p2 ^ 1'd1);

assign xor_ln895_79_fu_8574_p2 = (tmp_217_fu_8449_p3 ^ 1'd1);

assign xor_ln895_80_fu_9028_p2 = (tmp_223_fu_9012_p3 ^ 1'd1);

assign xor_ln895_81_fu_9078_p2 = (tmp_225_fu_9062_p3 ^ 1'd1);

assign xor_ln895_82_fu_9242_p2 = (xor_ln888_47_fu_9204_p2 ^ 1'd1);

assign xor_ln895_83_fu_9254_p2 = (tmp_227_fu_9129_p3 ^ 1'd1);

assign xor_ln895_84_fu_9521_p2 = (tmp_233_fu_9505_p3 ^ 1'd1);

assign xor_ln895_85_fu_2861_p2 = (xor_ln888_49_fu_2824_p2 ^ 1'd1);

assign xor_ln895_86_fu_2873_p2 = (tmp_235_fu_2745_p3 ^ 1'd1);

assign xor_ln895_87_fu_3614_p2 = (xor_ln888_51_fu_3582_p2 ^ 1'd1);

assign xor_ln895_88_fu_3626_p2 = (tmp_241_fu_3505_p3 ^ 1'd1);

assign xor_ln895_89_fu_4323_p2 = (tmp_247_fu_4307_p3 ^ 1'd1);

assign xor_ln895_90_fu_4373_p2 = (tmp_249_fu_4357_p3 ^ 1'd1);

assign xor_ln895_91_fu_4423_p2 = (tmp_251_fu_4407_p3 ^ 1'd1);

assign xor_ln895_92_fu_4473_p2 = (tmp_253_fu_4457_p3 ^ 1'd1);

assign xor_ln895_93_fu_5929_p2 = (xor_ln888_53_fu_5897_p2 ^ 1'd1);

assign xor_ln895_94_fu_5941_p2 = (tmp_255_fu_5820_p3 ^ 1'd1);

assign xor_ln895_95_fu_6614_p2 = (xor_ln888_55_fu_6576_p2 ^ 1'd1);

assign xor_ln895_96_fu_6626_p2 = (tmp_261_fu_6501_p3 ^ 1'd1);

assign xor_ln895_97_fu_7138_p2 = (tmp_267_fu_7122_p3 ^ 1'd1);

assign xor_ln895_98_fu_7188_p2 = (tmp_269_fu_7172_p3 ^ 1'd1);

assign xor_ln895_99_fu_7348_p2 = (xor_ln888_57_fu_7316_p2 ^ 1'd1);

assign xor_ln895_fu_1345_p2 = (tmp_fu_1323_p3 ^ 1'd1);

assign xor_ln896_100_fu_13333_p2 = (tmp_360_fu_13325_p3 ^ 1'd1);

assign xor_ln896_101_fu_13425_p2 = (1'd1 ^ and_ln890_40_fu_13389_p2);

assign xor_ln896_102_fu_7075_p2 = (or_ln896_20_fu_7069_p2 ^ and_ln891_20_fu_7033_p2);

assign xor_ln896_103_fu_7809_p2 = (or_ln896_21_fu_7803_p2 ^ and_ln891_21_fu_7767_p2);

assign xor_ln896_104_fu_13503_p2 = (tmp_370_fu_13495_p3 ^ 1'd1);

assign xor_ln896_105_fu_13595_p2 = (1'd1 ^ and_ln890_41_fu_13559_p2);

assign xor_ln896_106_fu_15239_p2 = (tmp_376_fu_15231_p3 ^ 1'd1);

assign xor_ln896_107_fu_15321_p2 = (1'd1 ^ and_ln890_42_fu_15291_p2);

assign xor_ln896_108_fu_8598_p2 = (or_ln896_22_fu_8592_p2 ^ and_ln891_22_fu_8556_p2);

assign xor_ln896_109_fu_13693_p2 = (tmp_384_fu_13685_p3 ^ 1'd1);

assign xor_ln896_10_fu_5354_p2 = (tmp_104_fu_5346_p3 ^ 1'd1);

assign xor_ln896_110_fu_13785_p2 = (1'd1 ^ and_ln890_43_fu_13749_p2);

assign xor_ln896_111_fu_15431_p2 = (tmp_390_fu_15423_p3 ^ 1'd1);

assign xor_ln896_112_fu_15513_p2 = (1'd1 ^ and_ln890_44_fu_15483_p2);

assign xor_ln896_113_fu_9278_p2 = (or_ln896_23_fu_9272_p2 ^ and_ln891_23_fu_9236_p2);

assign xor_ln896_114_fu_13867_p2 = (tmp_398_fu_13859_p3 ^ 1'd1);

assign xor_ln896_115_fu_13959_p2 = (1'd1 ^ and_ln890_45_fu_13923_p2);

assign xor_ln896_116_fu_15593_p2 = (tmp_404_fu_15585_p3 ^ 1'd1);

assign xor_ln896_117_fu_15687_p2 = (1'd1 ^ and_ln890_46_fu_15651_p2);

assign xor_ln896_118_fu_17379_p2 = (tmp_410_fu_17371_p3 ^ 1'd1);

assign xor_ln896_119_fu_17473_p2 = (1'd1 ^ and_ln890_47_fu_17437_p2);

assign xor_ln896_11_fu_5448_p2 = (1'd1 ^ and_ln890_5_fu_5412_p2);

assign xor_ln896_120_fu_14064_p2 = (tmp_416_fu_14056_p3 ^ 1'd1);

assign xor_ln896_121_fu_14156_p2 = (1'd1 ^ and_ln890_48_fu_14120_p2);

assign xor_ln896_122_fu_15830_p2 = (tmp_422_fu_15822_p3 ^ 1'd1);

assign xor_ln896_123_fu_15924_p2 = (1'd1 ^ and_ln890_49_fu_15888_p2);

assign xor_ln896_124_fu_17591_p2 = (tmp_428_fu_17583_p3 ^ 1'd1);

assign xor_ln896_125_fu_17685_p2 = (1'd1 ^ and_ln890_50_fu_17649_p2);

assign xor_ln896_126_fu_16025_p2 = (tmp_434_fu_16017_p3 ^ 1'd1);

assign xor_ln896_127_fu_16117_p2 = (1'd1 ^ and_ln890_51_fu_16081_p2);

assign xor_ln896_128_fu_2897_p2 = (or_ln896_24_fu_2891_p2 ^ and_ln891_24_fu_2855_p2);

assign xor_ln896_129_fu_4278_p2 = (or_ln896_25_reg_22626 ^ and_ln891_25_fu_4273_p2);

assign xor_ln896_12_fu_6044_p2 = (tmp_110_fu_6036_p3 ^ 1'd1);

assign xor_ln896_130_fu_16199_p2 = (tmp_444_fu_16191_p3 ^ 1'd1);

assign xor_ln896_131_fu_16291_p2 = (1'd1 ^ and_ln890_52_fu_16255_p2);

assign xor_ln896_132_fu_6442_p2 = (or_ln896_26_reg_22871 ^ and_ln891_26_fu_6437_p2);

assign xor_ln896_133_fu_6650_p2 = (or_ln896_27_fu_6644_p2 ^ and_ln891_27_fu_6608_p2);

assign xor_ln896_134_fu_14241_p2 = (tmp_454_fu_14233_p3 ^ 1'd1);

assign xor_ln896_135_fu_14333_p2 = (1'd1 ^ and_ln890_53_fu_14297_p2);

assign xor_ln896_136_fu_16397_p2 = (tmp_460_fu_16389_p3 ^ 1'd1);

assign xor_ln896_137_fu_16479_p2 = (1'd1 ^ and_ln890_54_fu_16449_p2);

assign xor_ln896_138_fu_7843_p2 = (or_ln896_28_reg_22998 ^ and_ln891_28_fu_7838_p2);

assign xor_ln896_139_fu_14431_p2 = (tmp_468_fu_14423_p3 ^ 1'd1);

assign xor_ln896_13_fu_6138_p2 = (1'd1 ^ and_ln890_6_fu_6102_p2);

assign xor_ln896_140_fu_14523_p2 = (1'd1 ^ and_ln890_55_fu_14487_p2);

assign xor_ln896_141_fu_16589_p2 = (tmp_474_fu_16581_p3 ^ 1'd1);

assign xor_ln896_142_fu_16671_p2 = (1'd1 ^ and_ln890_56_fu_16641_p2);

assign xor_ln896_143_fu_8625_p2 = (or_ln896_29_reg_23064 ^ and_ln891_29_fu_8620_p2);

assign xor_ln896_144_fu_14605_p2 = (tmp_482_fu_14597_p3 ^ 1'd1);

assign xor_ln896_145_fu_14697_p2 = (1'd1 ^ and_ln890_57_fu_14661_p2);

assign xor_ln896_146_fu_16751_p2 = (tmp_488_fu_16743_p3 ^ 1'd1);

assign xor_ln896_147_fu_16845_p2 = (1'd1 ^ and_ln890_58_fu_16809_p2);

assign xor_ln896_148_fu_18207_p2 = (tmp_494_fu_18199_p3 ^ 1'd1);

assign xor_ln896_149_fu_18301_p2 = (1'd1 ^ and_ln890_59_fu_18265_p2);

assign xor_ln896_14_fu_6740_p2 = (tmp_116_fu_6732_p3 ^ 1'd1);

assign xor_ln896_150_fu_14802_p2 = (tmp_500_fu_14794_p3 ^ 1'd1);

assign xor_ln896_151_fu_14894_p2 = (1'd1 ^ and_ln890_60_fu_14858_p2);

assign xor_ln896_152_fu_16988_p2 = (tmp_506_fu_16980_p3 ^ 1'd1);

assign xor_ln896_153_fu_17082_p2 = (1'd1 ^ and_ln890_61_fu_17046_p2);

assign xor_ln896_154_fu_18419_p2 = (tmp_512_fu_18411_p3 ^ 1'd1);

assign xor_ln896_155_fu_18513_p2 = (1'd1 ^ and_ln890_62_fu_18477_p2);

assign xor_ln896_156_fu_10522_p2 = (or_ln896_30_fu_10516_p2 ^ and_ln891_30_fu_10480_p2);

assign xor_ln896_157_fu_11085_p2 = (or_ln896_31_fu_11079_p2 ^ and_ln891_31_fu_11043_p2);

assign xor_ln896_158_fu_11760_p2 = (or_ln896_32_fu_11754_p2 ^ and_ln891_32_fu_11718_p2);

assign xor_ln896_159_fu_12439_p2 = (1'd1 ^ and_ln896_63_fu_12433_p2);

assign xor_ln896_15_fu_6834_p2 = (1'd1 ^ and_ln890_7_fu_6798_p2);

assign xor_ln896_160_fu_10712_p2 = (or_ln896_33_fu_10706_p2 ^ and_ln891_33_fu_10670_p2);

assign xor_ln896_161_fu_12596_p2 = (1'd1 ^ and_ln896_65_fu_12590_p2);

assign xor_ln896_162_fu_11315_p2 = (or_ln896_34_fu_11309_p2 ^ and_ln891_34_fu_11273_p2);

assign xor_ln896_163_fu_11956_p2 = (or_ln896_35_fu_11950_p2 ^ and_ln891_35_fu_11914_p2);

assign xor_ln896_164_fu_10886_p2 = (or_ln896_36_fu_10880_p2 ^ and_ln891_36_fu_10844_p2);

assign xor_ln896_165_fu_11564_p2 = (or_ln896_37_fu_11558_p2 ^ and_ln891_37_fu_11522_p2);

assign xor_ln896_166_fu_12162_p2 = (or_ln896_38_fu_12156_p2 ^ and_ln891_38_fu_12120_p2);

assign xor_ln896_167_fu_13263_p2 = (or_ln896_39_fu_13257_p2 ^ and_ln891_39_fu_13221_p2);

assign xor_ln896_168_fu_13437_p2 = (or_ln896_40_fu_13431_p2 ^ and_ln891_40_fu_13395_p2);

assign xor_ln896_169_fu_13607_p2 = (or_ln896_41_fu_13601_p2 ^ and_ln891_41_fu_13565_p2);

assign xor_ln896_16_fu_7452_p2 = (tmp_122_fu_7444_p3 ^ 1'd1);

assign xor_ln896_170_fu_17144_p2 = (or_ln896_42_reg_23635 ^ and_ln891_42_fu_17139_p2);

assign xor_ln896_171_fu_13797_p2 = (or_ln896_43_fu_13791_p2 ^ and_ln891_43_fu_13755_p2);

assign xor_ln896_172_fu_17232_p2 = (or_ln896_44_reg_23671 ^ and_ln891_44_fu_17227_p2);

assign xor_ln896_173_fu_13971_p2 = (or_ln896_45_fu_13965_p2 ^ and_ln891_45_fu_13929_p2);

assign xor_ln896_174_fu_15699_p2 = (or_ln896_46_fu_15693_p2 ^ and_ln891_46_fu_15657_p2);

assign xor_ln896_175_fu_17485_p2 = (or_ln896_47_fu_17479_p2 ^ and_ln891_47_fu_17443_p2);

assign xor_ln896_176_fu_14168_p2 = (or_ln896_48_fu_14162_p2 ^ and_ln891_48_fu_14126_p2);

assign xor_ln896_177_fu_15936_p2 = (or_ln896_49_fu_15930_p2 ^ and_ln891_49_fu_15894_p2);

assign xor_ln896_178_fu_17697_p2 = (or_ln896_50_fu_17691_p2 ^ and_ln891_50_fu_17655_p2);

assign xor_ln896_179_fu_16129_p2 = (or_ln896_51_fu_16123_p2 ^ and_ln891_51_fu_16087_p2);

assign xor_ln896_17_fu_7546_p2 = (1'd1 ^ and_ln890_8_fu_7510_p2);

assign xor_ln896_180_fu_16303_p2 = (or_ln896_52_fu_16297_p2 ^ and_ln891_52_fu_16261_p2);

assign xor_ln896_181_fu_14345_p2 = (or_ln896_53_fu_14339_p2 ^ and_ln891_53_fu_14303_p2);

assign xor_ln896_182_fu_17972_p2 = (or_ln896_54_reg_23769 ^ and_ln891_54_fu_17967_p2);

assign xor_ln896_183_fu_14535_p2 = (or_ln896_55_fu_14529_p2 ^ and_ln891_55_fu_14493_p2);

assign xor_ln896_184_fu_18060_p2 = (or_ln896_56_reg_23805 ^ and_ln891_56_fu_18055_p2);

assign xor_ln896_185_fu_14709_p2 = (or_ln896_57_fu_14703_p2 ^ and_ln891_57_fu_14667_p2);

assign xor_ln896_186_fu_16857_p2 = (or_ln896_58_fu_16851_p2 ^ and_ln891_58_fu_16815_p2);

assign xor_ln896_187_fu_18313_p2 = (or_ln896_59_fu_18307_p2 ^ and_ln891_59_fu_18271_p2);

assign xor_ln896_188_fu_14906_p2 = (or_ln896_60_fu_14900_p2 ^ and_ln891_60_fu_14864_p2);

assign xor_ln896_189_fu_17094_p2 = (or_ln896_61_fu_17088_p2 ^ and_ln891_61_fu_17052_p2);

assign xor_ln896_18_fu_8245_p2 = (tmp_128_fu_8237_p3 ^ 1'd1);

assign xor_ln896_190_fu_18525_p2 = (or_ln896_62_fu_18519_p2 ^ and_ln891_62_fu_18483_p2);

assign xor_ln896_191_fu_12706_p2 = (1'd1 ^ and_ln896_67_fu_12700_p2);

assign xor_ln896_192_fu_12927_p2 = (1'd1 ^ and_ln896_69_fu_12921_p2);

assign xor_ln896_193_fu_13076_p2 = (1'd1 ^ and_ln896_71_fu_13070_p2);

assign xor_ln896_19_fu_8339_p2 = (1'd1 ^ and_ln890_9_fu_8303_p2);

assign xor_ln896_1_fu_2117_p2 = (1'd1 ^ and_ln890_fu_2081_p2);

assign xor_ln896_20_fu_8859_p2 = (tmp_134_fu_8851_p3 ^ 1'd1);

assign xor_ln896_21_fu_8953_p2 = (1'd1 ^ and_ln890_10_fu_8917_p2);

assign xor_ln896_22_fu_9368_p2 = (tmp_140_fu_9360_p3 ^ 1'd1);

assign xor_ln896_23_fu_9462_p2 = (1'd1 ^ and_ln890_11_fu_9426_p2);

assign xor_ln896_24_fu_9729_p2 = (tmp_146_fu_9721_p3 ^ 1'd1);

assign xor_ln896_25_fu_9823_p2 = (1'd1 ^ and_ln890_12_fu_9787_p2);

assign xor_ln896_26_fu_2129_p2 = (or_ln896_fu_2123_p2 ^ and_ln891_fu_2087_p2);

assign xor_ln896_27_fu_2496_p2 = (or_ln896_1_fu_2490_p2 ^ and_ln891_1_fu_2454_p2);

assign xor_ln896_28_fu_10040_p2 = (tmp_156_fu_10032_p3 ^ 1'd1);

assign xor_ln896_29_fu_10134_p2 = (1'd1 ^ and_ln890_13_fu_10098_p2);

assign xor_ln896_2_fu_2390_p2 = (tmp_80_fu_2382_p3 ^ 1'd1);

assign xor_ln896_30_fu_3245_p2 = (or_ln896_2_fu_3239_p2 ^ and_ln891_2_fu_3203_p2);

assign xor_ln896_31_fu_3998_p2 = (or_ln896_3_fu_3992_p2 ^ and_ln891_3_fu_3956_p2);

assign xor_ln896_32_fu_2600_p2 = (tmp_166_fu_2592_p3 ^ 1'd1);

assign xor_ln896_33_fu_2692_p2 = (1'd1 ^ and_ln890_14_fu_2656_p2);

assign xor_ln896_34_fu_3382_p2 = (tmp_172_fu_3374_p3 ^ 1'd1);

assign xor_ln896_35_fu_3464_p2 = (1'd1 ^ and_ln890_15_fu_3434_p2);

assign xor_ln896_36_fu_4141_p2 = (tmp_178_fu_4133_p3 ^ 1'd1);

assign xor_ln896_37_fu_4235_p2 = (1'd1 ^ and_ln890_16_fu_4199_p2);

assign xor_ln896_38_fu_5000_p2 = (tmp_184_fu_4992_p3 ^ 1'd1);

assign xor_ln896_39_fu_5094_p2 = (1'd1 ^ and_ln890_17_fu_5058_p2);

assign xor_ln896_3_fu_2484_p2 = (1'd1 ^ and_ln890_1_fu_2448_p2);

assign xor_ln896_40_fu_4839_p2 = (or_ln896_4_fu_4833_p2 ^ and_ln891_4_fu_4797_p2);

assign xor_ln896_41_fu_5460_p2 = (or_ln896_5_fu_5454_p2 ^ and_ln891_5_fu_5418_p2);

assign xor_ln896_42_fu_5690_p2 = (tmp_194_fu_5682_p3 ^ 1'd1);

assign xor_ln896_43_fu_5772_p2 = (1'd1 ^ and_ln890_18_fu_5742_p2);

assign xor_ln896_44_fu_6302_p2 = (tmp_200_fu_6294_p3 ^ 1'd1);

assign xor_ln896_45_fu_6396_p2 = (1'd1 ^ and_ln890_19_fu_6360_p2);

assign xor_ln896_46_fu_6969_p2 = (tmp_206_fu_6961_p3 ^ 1'd1);

assign xor_ln896_47_fu_7063_p2 = (1'd1 ^ and_ln890_20_fu_7027_p2);

assign xor_ln896_48_fu_7703_p2 = (tmp_212_fu_7695_p3 ^ 1'd1);

assign xor_ln896_49_fu_7797_p2 = (1'd1 ^ and_ln890_21_fu_7761_p2);

assign xor_ln896_4_fu_3139_p2 = (tmp_86_fu_3131_p3 ^ 1'd1);

assign xor_ln896_50_fu_6150_p2 = (or_ln896_6_fu_6144_p2 ^ and_ln891_6_fu_6108_p2);

assign xor_ln896_51_fu_8492_p2 = (tmp_220_fu_8484_p3 ^ 1'd1);

assign xor_ln896_52_fu_8586_p2 = (1'd1 ^ and_ln890_22_fu_8550_p2);

assign xor_ln896_53_fu_6846_p2 = (or_ln896_7_fu_6840_p2 ^ and_ln891_7_fu_6804_p2);

assign xor_ln896_54_fu_7558_p2 = (or_ln896_8_fu_7552_p2 ^ and_ln891_8_fu_7516_p2);

assign xor_ln896_55_fu_9172_p2 = (tmp_230_fu_9164_p3 ^ 1'd1);

assign xor_ln896_56_fu_9266_p2 = (1'd1 ^ and_ln890_23_fu_9230_p2);

assign xor_ln896_57_fu_8351_p2 = (or_ln896_9_fu_8345_p2 ^ and_ln891_9_fu_8309_p2);

assign xor_ln896_58_fu_2793_p2 = (tmp_238_fu_2785_p3 ^ 1'd1);

assign xor_ln896_59_fu_2885_p2 = (1'd1 ^ and_ln890_24_fu_2849_p2);

assign xor_ln896_5_fu_3233_p2 = (1'd1 ^ and_ln890_2_fu_3197_p2);

assign xor_ln896_60_fu_3556_p2 = (tmp_244_fu_3548_p3 ^ 1'd1);

assign xor_ln896_61_fu_3638_p2 = (1'd1 ^ and_ln890_25_fu_3608_p2);

assign xor_ln896_62_fu_8965_p2 = (or_ln896_10_fu_8959_p2 ^ and_ln891_10_fu_8923_p2);

assign xor_ln896_63_fu_9474_p2 = (or_ln896_11_fu_9468_p2 ^ and_ln891_11_fu_9432_p2);

assign xor_ln896_64_fu_9835_p2 = (or_ln896_12_fu_9829_p2 ^ and_ln891_12_fu_9793_p2);

assign xor_ln896_65_fu_10146_p2 = (or_ln896_13_fu_10140_p2 ^ and_ln891_13_fu_10104_p2);

assign xor_ln896_66_fu_5871_p2 = (tmp_258_fu_5863_p3 ^ 1'd1);

assign xor_ln896_67_fu_5953_p2 = (1'd1 ^ and_ln890_26_fu_5923_p2);

assign xor_ln896_68_fu_6544_p2 = (tmp_264_fu_6536_p3 ^ 1'd1);

assign xor_ln896_69_fu_6638_p2 = (1'd1 ^ and_ln890_27_fu_6602_p2);

assign xor_ln896_6_fu_3892_p2 = (tmp_92_fu_3884_p3 ^ 1'd1);

assign xor_ln896_70_fu_2704_p2 = (or_ln896_14_fu_2698_p2 ^ and_ln891_14_fu_2662_p2);

assign xor_ln896_71_fu_4043_p2 = (or_ln896_15_reg_22590 ^ and_ln891_15_fu_4038_p2);

assign xor_ln896_72_fu_7290_p2 = (tmp_274_fu_7282_p3 ^ 1'd1);

assign xor_ln896_73_fu_7372_p2 = (1'd1 ^ and_ln890_28_fu_7342_p2);

assign xor_ln896_74_fu_4247_p2 = (or_ln896_16_fu_4241_p2 ^ and_ln891_16_fu_4205_p2);

assign xor_ln896_75_fu_5106_p2 = (or_ln896_17_fu_5100_p2 ^ and_ln891_17_fu_5064_p2);

assign xor_ln896_76_fu_8040_p2 = (tmp_284_fu_8032_p3 ^ 1'd1);

assign xor_ln896_77_fu_8122_p2 = (1'd1 ^ and_ln890_29_fu_8092_p2);

assign xor_ln896_78_fu_10418_p2 = (tmp_296_fu_10410_p3 ^ 1'd1);

assign xor_ln896_79_fu_10510_p2 = (1'd1 ^ and_ln890_30_fu_10474_p2);

assign xor_ln896_7_fu_3986_p2 = (1'd1 ^ and_ln890_3_fu_3950_p2);

assign xor_ln896_80_fu_10979_p2 = (tmp_302_fu_10971_p3 ^ 1'd1);

assign xor_ln896_81_fu_11073_p2 = (1'd1 ^ and_ln890_31_fu_11037_p2);

assign xor_ln896_82_fu_11654_p2 = (tmp_308_fu_11646_p3 ^ 1'd1);

assign xor_ln896_83_fu_11748_p2 = (1'd1 ^ and_ln890_32_fu_11712_p2);

assign xor_ln896_84_fu_10608_p2 = (tmp_314_fu_10600_p3 ^ 1'd1);

assign xor_ln896_85_fu_10700_p2 = (1'd1 ^ and_ln890_33_fu_10664_p2);

assign xor_ln896_86_fu_11209_p2 = (tmp_320_fu_11201_p3 ^ 1'd1);

assign xor_ln896_87_fu_11303_p2 = (1'd1 ^ and_ln890_34_fu_11267_p2);

assign xor_ln896_88_fu_11850_p2 = (tmp_326_fu_11842_p3 ^ 1'd1);

assign xor_ln896_89_fu_11944_p2 = (1'd1 ^ and_ln890_35_fu_11908_p2);

assign xor_ln896_8_fu_4733_p2 = (tmp_98_fu_4725_p3 ^ 1'd1);

assign xor_ln896_90_fu_10782_p2 = (tmp_332_fu_10774_p3 ^ 1'd1);

assign xor_ln896_91_fu_10874_p2 = (1'd1 ^ and_ln890_36_fu_10838_p2);

assign xor_ln896_92_fu_11458_p2 = (tmp_338_fu_11450_p3 ^ 1'd1);

assign xor_ln896_93_fu_11552_p2 = (1'd1 ^ and_ln890_37_fu_11516_p2);

assign xor_ln896_94_fu_12056_p2 = (tmp_344_fu_12048_p3 ^ 1'd1);

assign xor_ln896_95_fu_12150_p2 = (1'd1 ^ and_ln890_38_fu_12114_p2);

assign xor_ln896_96_fu_13159_p2 = (tmp_350_fu_13151_p3 ^ 1'd1);

assign xor_ln896_97_fu_13251_p2 = (1'd1 ^ and_ln890_39_fu_13215_p2);

assign xor_ln896_98_fu_6200_p2 = (or_ln896_18_reg_22819 ^ and_ln891_18_fu_6195_p2);

assign xor_ln896_99_fu_6408_p2 = (or_ln896_19_fu_6402_p2 ^ and_ln891_19_fu_6366_p2);

assign xor_ln896_9_fu_4827_p2 = (1'd1 ^ and_ln890_4_fu_4791_p2);

assign xor_ln896_fu_2025_p2 = (tmp_74_fu_2017_p3 ^ 1'd1);

assign zext_ln377_10_fu_8842_p1 = tmp_133_reg_22772;

assign zext_ln377_11_fu_9351_p1 = tmp_139_reg_22783;

assign zext_ln377_12_fu_9712_p1 = tmp_145_reg_22902;

assign zext_ln377_13_fu_10023_p1 = tmp_155_reg_22957;

assign zext_ln377_14_fu_2582_p1 = tmp_165_fu_2575_p3;

assign zext_ln377_15_fu_3364_p1 = tmp_171_fu_3357_p3;

assign zext_ln377_16_fu_4124_p1 = tmp_177_reg_22506;

assign zext_ln377_17_fu_4983_p1 = tmp_183_reg_22420;

assign zext_ln377_18_fu_5673_p1 = tmp_193_reg_22740;

assign zext_ln377_19_fu_6285_p1 = tmp_199_reg_22751;

assign zext_ln377_1_fu_2373_p1 = tmp_79_reg_22436;

assign zext_ln377_20_fu_6952_p1 = tmp_205_reg_22830;

assign zext_ln377_21_fu_7685_p1 = tmp_211_fu_7677_p3;

assign zext_ln377_22_fu_8475_p1 = tmp_219_reg_22927;

assign zext_ln377_23_fu_9155_p1 = tmp_229_reg_23028;

assign zext_ln377_24_fu_2775_p1 = tmp_237_fu_2768_p3;

assign zext_ln377_25_fu_3538_p1 = tmp_243_fu_3531_p3;

assign zext_ln377_26_fu_5853_p1 = tmp_257_fu_5846_p3;

assign zext_ln377_27_fu_6527_p1 = tmp_263_reg_22882;

assign zext_ln377_28_fu_7272_p1 = tmp_273_fu_7265_p3;

assign zext_ln377_29_fu_8022_p1 = tmp_283_fu_8015_p3;

assign zext_ln377_2_fu_3122_p1 = tmp_85_reg_22468;

assign zext_ln377_30_fu_10400_p1 = tmp_295_fu_10393_p3;

assign zext_ln377_31_fu_10962_p1 = tmp_301_reg_23249;

assign zext_ln377_32_fu_11637_p1 = tmp_307_reg_23197;

assign zext_ln377_33_fu_10590_p1 = tmp_313_fu_10583_p3;

assign zext_ln377_34_fu_11192_p1 = tmp_319_reg_23260;

assign zext_ln377_35_fu_11833_p1 = tmp_325_reg_23115;

assign zext_ln377_36_fu_10764_p1 = tmp_331_fu_10757_p3;

assign zext_ln377_37_fu_11441_p1 = tmp_337_reg_23171;

assign zext_ln377_38_fu_12039_p1 = tmp_343_reg_23208;

assign zext_ln377_39_fu_13141_p1 = tmp_349_fu_13134_p3;

assign zext_ln377_3_fu_3875_p1 = tmp_91_reg_22405;

assign zext_ln377_40_fu_13315_p1 = tmp_359_fu_13308_p3;

assign zext_ln377_41_fu_13485_p1 = tmp_369_fu_13478_p3;

assign zext_ln377_42_fu_15221_p1 = tmp_375_fu_15214_p3;

assign zext_ln377_43_fu_13675_p1 = tmp_383_fu_13668_p3;

assign zext_ln377_44_fu_15413_p1 = tmp_389_fu_15406_p3;

assign zext_ln377_45_fu_13849_p1 = tmp_397_fu_13842_p3;

assign zext_ln377_46_fu_15576_p1 = tmp_403_reg_23511;

assign zext_ln377_47_fu_17362_p1 = tmp_409_reg_23687;

assign zext_ln377_48_fu_14046_p1 = tmp_415_fu_14039_p3;

assign zext_ln377_49_fu_15813_p1 = tmp_421_reg_23537;

assign zext_ln377_4_fu_4716_p1 = tmp_97_reg_22479;

assign zext_ln377_50_fu_17574_p1 = tmp_427_reg_23703;

assign zext_ln377_51_fu_16007_p1 = tmp_433_fu_16000_p3;

assign zext_ln377_52_fu_16181_p1 = tmp_443_fu_16174_p3;

assign zext_ln377_53_fu_14223_p1 = tmp_453_fu_14216_p3;

assign zext_ln377_54_fu_16379_p1 = tmp_459_fu_16372_p3;

assign zext_ln377_55_fu_14413_p1 = tmp_467_fu_14406_p3;

assign zext_ln377_56_fu_16571_p1 = tmp_473_fu_16564_p3;

assign zext_ln377_57_fu_14587_p1 = tmp_481_fu_14580_p3;

assign zext_ln377_58_fu_16734_p1 = tmp_487_reg_23573;

assign zext_ln377_59_fu_18190_p1 = tmp_493_reg_23821;

assign zext_ln377_5_fu_5337_p1 = tmp_103_reg_22533;

assign zext_ln377_60_fu_14784_p1 = tmp_499_fu_14777_p3;

assign zext_ln377_61_fu_16971_p1 = tmp_505_reg_23599;

assign zext_ln377_62_fu_18402_p1 = tmp_511_reg_23837;

assign zext_ln377_6_fu_6027_p1 = tmp_109_reg_22652;

assign zext_ln377_7_fu_6723_p1 = tmp_115_reg_22663;

assign zext_ln377_8_fu_7435_p1 = tmp_121_reg_22709;

assign zext_ln377_9_fu_8227_p1 = tmp_127_fu_8219_p3;

assign zext_ln377_fu_2007_p1 = tmp_73_fu_2000_p3;

assign zext_ln50_10_fu_19593_p1 = select_ln49_10_fu_19585_p3;

assign zext_ln50_11_fu_19610_p1 = select_ln49_11_fu_19602_p3;

assign zext_ln50_12_fu_19769_p1 = select_ln49_12_fu_19761_p3;

assign zext_ln50_13_fu_19786_p1 = select_ln49_13_fu_19778_p3;

assign zext_ln50_14_fu_19945_p1 = select_ln49_14_fu_19937_p3;

assign zext_ln50_15_fu_19962_p1 = select_ln49_15_fu_19954_p3;

assign zext_ln50_16_fu_20121_p1 = select_ln49_16_fu_20113_p3;

assign zext_ln50_17_fu_20138_p1 = select_ln49_17_fu_20130_p3;

assign zext_ln50_1_fu_18730_p1 = select_ln49_1_fu_18722_p3;

assign zext_ln50_2_fu_18889_p1 = select_ln49_2_fu_18881_p3;

assign zext_ln50_3_fu_18906_p1 = select_ln49_3_fu_18898_p3;

assign zext_ln50_4_fu_19065_p1 = select_ln49_4_fu_19057_p3;

assign zext_ln50_5_fu_19082_p1 = select_ln49_5_fu_19074_p3;

assign zext_ln50_6_fu_19241_p1 = select_ln49_6_fu_19233_p3;

assign zext_ln50_7_fu_19258_p1 = select_ln49_7_fu_19250_p3;

assign zext_ln50_8_fu_19417_p1 = select_ln49_8_fu_19409_p3;

assign zext_ln50_9_fu_19434_p1 = select_ln49_9_fu_19426_p3;

assign zext_ln50_fu_18713_p1 = select_ln49_fu_18705_p3;

endmodule //mpc_qp_admm
